<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-81.8804,90.472,173.486,-38.6125</PageViewport>
<gate>
<ID>780</ID>
<type>DE_TO</type>
<position>13,32.5</position>
<input>
<ID>IN_0</ID>522 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID USE-USER-INSTRUCTION</lparam></gate>
<gate>
<ID>392</ID>
<type>AE_REGISTER8</type>
<position>33,56.5</position>
<input>
<ID>IN_0</ID>437 </input>
<input>
<ID>IN_1</ID>449 </input>
<input>
<ID>IN_2</ID>463 </input>
<input>
<ID>IN_3</ID>481 </input>
<input>
<ID>IN_4</ID>515 </input>
<input>
<ID>IN_5</ID>405 </input>
<input>
<ID>IN_6</ID>383 </input>
<input>
<ID>IN_7</ID>382 </input>
<output>
<ID>OUT_0</ID>287 </output>
<output>
<ID>OUT_1</ID>288 </output>
<output>
<ID>OUT_2</ID>384 </output>
<output>
<ID>OUT_3</ID>385 </output>
<output>
<ID>OUT_4</ID>291 </output>
<output>
<ID>OUT_5</ID>292 </output>
<output>
<ID>OUT_6</ID>293 </output>
<output>
<ID>OUT_7</ID>294 </output>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>load</ID>358 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 106</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>394</ID>
<type>DE_TO</type>
<position>41.5,48</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-0</lparam></gate>
<gate>
<ID>395</ID>
<type>DE_TO</type>
<position>41.5,65.5</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-REG</lparam></gate>
<gate>
<ID>396</ID>
<type>DE_TO</type>
<position>41.5,63</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-3</lparam></gate>
<gate>
<ID>397</ID>
<type>DE_TO</type>
<position>41.5,60.5</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-2</lparam></gate>
<gate>
<ID>398</ID>
<type>DE_TO</type>
<position>41.5,58</position>
<input>
<ID>IN_0</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-1</lparam></gate>
<gate>
<ID>399</ID>
<type>DE_TO</type>
<position>41.5,55.5</position>
<input>
<ID>IN_0</ID>385 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-0</lparam></gate>
<gate>
<ID>400</ID>
<type>DE_TO</type>
<position>41.5,53</position>
<input>
<ID>IN_0</ID>384 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-2</lparam></gate>
<gate>
<ID>790</ID>
<type>DE_TO</type>
<position>13,30</position>
<input>
<ID>IN_0</ID>663 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WRITE-INSTRUCTION</lparam></gate>
<gate>
<ID>401</ID>
<type>DE_TO</type>
<position>41.5,50.5</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_REGISTER4</type>
<position>-19.5,-13</position>
<output>
<ID>OUT_0</ID>24 </output>
<output>
<ID>OUT_1</ID>23 </output>
<output>
<ID>OUT_2</ID>22 </output>
<output>
<ID>OUT_3</ID>21 </output>
<input>
<ID>clear</ID>583 </input>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>count_enable</ID>51 </input>
<input>
<ID>count_up</ID>51 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>17</ID>
<type>EE_VDD</type>
<position>-6.5,64.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>796</ID>
<type>DD_KEYPAD_HEX</type>
<position>13,19</position>
<output>
<ID>OUT_0</ID>81 </output>
<output>
<ID>OUT_1</ID>83 </output>
<output>
<ID>OUT_2</ID>82 </output>
<output>
<ID>OUT_3</ID>80 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>407</ID>
<type>AA_LABEL</type>
<position>35.5,67.5</position>
<gparam>LABEL_TEXT IR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_REGISTER4</type>
<position>43,-5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>9 </input>
<output>
<ID>OUT_0</ID>15 </output>
<output>
<ID>OUT_1</ID>16 </output>
<output>
<ID>OUT_2</ID>17 </output>
<output>
<ID>OUT_3</ID>14 </output>
<input>
<ID>clear</ID>154 </input>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>load</ID>141 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 13</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>408</ID>
<type>DE_TO</type>
<position>-3,60</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-3</lparam></gate>
<gate>
<ID>409</ID>
<type>DE_TO</type>
<position>-3,57.5</position>
<input>
<ID>IN_0</ID>307 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>43.5,5.5</position>
<gparam>LABEL_TEXT MAR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>410</ID>
<type>DE_TO</type>
<position>-3,55</position>
<input>
<ID>IN_0</ID>306 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-1</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>35.5,-1</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-3</lparam></gate>
<gate>
<ID>800</ID>
<type>DE_TO</type>
<position>-29,36</position>
<input>
<ID>IN_0</ID>627 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RUN-PROGRAM</lparam></gate>
<gate>
<ID>411</ID>
<type>DE_TO</type>
<position>-3,52.5</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-0</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>35.5,-8.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-0</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>35.5,-6</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-1</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>35.5,-3.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-2</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>51,-1</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-3</lparam></gate>
<gate>
<ID>804</ID>
<type>DE_TO</type>
<position>20,22</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-USER-3</lparam></gate>
<gate>
<ID>26</ID>
<type>DE_TO</type>
<position>51,-3.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-2</lparam></gate>
<gate>
<ID>805</ID>
<type>DE_TO</type>
<position>20,20</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-USER-2</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>51,-6</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-1</lparam></gate>
<gate>
<ID>806</ID>
<type>DE_TO</type>
<position>20,18</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-USER-1</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>-18,60</position>
<input>
<ID>IN_0</ID>317 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-3</lparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>51,-8.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-0</lparam></gate>
<gate>
<ID>807</ID>
<type>DE_TO</type>
<position>20,16</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-USER-0</lparam></gate>
<gate>
<ID>418</ID>
<type>DA_FROM</type>
<position>-18,52.5</position>
<input>
<ID>IN_0</ID>314 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-0</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_REGISTER4</type>
<position>82.5,-6</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<input>
<ID>IN_2</ID>139 </input>
<input>
<ID>IN_3</ID>140 </input>
<output>
<ID>OUT_0</ID>143 </output>
<output>
<ID>OUT_1</ID>144 </output>
<output>
<ID>OUT_2</ID>145 </output>
<input>
<ID>clear</ID>163 </input>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>load</ID>150 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>419</ID>
<type>DA_FROM</type>
<position>-18,55</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-33,41</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>809</ID>
<type>AA_LABEL</type>
<position>19.5,26.5</position>
<gparam>LABEL_TEXT Instruction Location</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>420</ID>
<type>DA_FROM</type>
<position>-18,57.5</position>
<input>
<ID>IN_0</ID>316 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-2</lparam></gate>
<gate>
<ID>31</ID>
<type>DE_TO</type>
<position>-29,41</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RESET-PC</lparam></gate>
<gate>
<ID>421</ID>
<type>AE_REGISTER8</type>
<position>79.5,55.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>310 </input>
<input>
<ID>IN_2</ID>311 </input>
<input>
<ID>IN_3</ID>312 </input>
<input>
<ID>IN_4</ID>313 </input>
<input>
<ID>IN_5</ID>326 </input>
<input>
<ID>IN_6</ID>327 </input>
<input>
<ID>IN_7</ID>304 </input>
<output>
<ID>OUT_0</ID>318 </output>
<output>
<ID>OUT_1</ID>319 </output>
<output>
<ID>OUT_2</ID>320 </output>
<output>
<ID>OUT_3</ID>321 </output>
<output>
<ID>OUT_4</ID>322 </output>
<output>
<ID>OUT_5</ID>323 </output>
<output>
<ID>OUT_6</ID>324 </output>
<output>
<ID>OUT_7</ID>325 </output>
<input>
<ID>clear</ID>553 </input>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>load</ID>359 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>422</ID>
<type>DE_TO</type>
<position>89,47.5</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-0</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>76,-8</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-0</lparam></gate>
<gate>
<ID>812</ID>
<type>AA_TOGGLE</type>
<position>-33,36</position>
<output>
<ID>OUT_0</ID>627 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>423</ID>
<type>DE_TO</type>
<position>89,65</position>
<input>
<ID>IN_0</ID>325 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-7</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>76,-6</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-1</lparam></gate>
<gate>
<ID>813</ID>
<type>AA_LABEL</type>
<position>-6.5,34</position>
<gparam>LABEL_TEXT IR Inputs</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>424</ID>
<type>DE_TO</type>
<position>89,62.5</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-6</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>76,-4</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-2</lparam></gate>
<gate>
<ID>425</ID>
<type>DE_TO</type>
<position>89,60</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-5</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>-15,-20</position>
<input>
<ID>IN_0</ID>583 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID SEQ-RESET</lparam></gate>
<gate>
<ID>426</ID>
<type>DE_TO</type>
<position>89,57.5</position>
<input>
<ID>IN_0</ID>322 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-4</lparam></gate>
<gate>
<ID>37</ID>
<type>BI_DECODER_4x16</type>
<position>-11.5,-6.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>22 </input>
<input>
<ID>IN_3</ID>21 </input>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>26 </output>
<output>
<ID>OUT_2</ID>27 </output>
<output>
<ID>OUT_3</ID>28 </output>
<output>
<ID>OUT_4</ID>29 </output>
<output>
<ID>OUT_5</ID>30 </output>
<output>
<ID>OUT_6</ID>31 </output>
<output>
<ID>OUT_7</ID>33 </output>
<output>
<ID>OUT_8</ID>34 </output>
<output>
<ID>OUT_9</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>427</ID>
<type>DE_TO</type>
<position>89,55</position>
<input>
<ID>IN_0</ID>321 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-3</lparam></gate>
<gate>
<ID>428</ID>
<type>DE_TO</type>
<position>89,52.5</position>
<input>
<ID>IN_0</ID>320 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-2</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>-3,-15.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-FETCH-2</lparam></gate>
<gate>
<ID>429</ID>
<type>DE_TO</type>
<position>89,50</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-1</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>-3,-17.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-FETCH-1</lparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>-3,-13.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-DECODE</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>-3,-11.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-1</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>-3,-9.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-2</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>-3,-7.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-3</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>-3,-5.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-4</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>-3,-3.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-5</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>-3,-1.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-6</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>-3,0.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-7</lparam></gate>
<gate>
<ID>438</ID>
<type>AE_REGISTER8</type>
<position>120.5,55.5</position>
<input>
<ID>IN_0</ID>284 </input>
<input>
<ID>IN_1</ID>267 </input>
<input>
<ID>IN_2</ID>332 </input>
<input>
<ID>IN_3</ID>333 </input>
<input>
<ID>IN_4</ID>342 </input>
<input>
<ID>IN_5</ID>343 </input>
<input>
<ID>IN_6</ID>330 </input>
<input>
<ID>IN_7</ID>329 </input>
<output>
<ID>OUT_0</ID>334 </output>
<output>
<ID>OUT_1</ID>335 </output>
<output>
<ID>OUT_2</ID>336 </output>
<output>
<ID>OUT_3</ID>337 </output>
<output>
<ID>OUT_4</ID>338 </output>
<output>
<ID>OUT_5</ID>339 </output>
<output>
<ID>OUT_6</ID>340 </output>
<output>
<ID>OUT_7</ID>341 </output>
<input>
<ID>clear</ID>554 </input>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>load</ID>360 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>439</ID>
<type>DE_TO</type>
<position>130,47.5</position>
<input>
<ID>IN_0</ID>334 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-0</lparam></gate>
<gate>
<ID>440</ID>
<type>DE_TO</type>
<position>130,65</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-7</lparam></gate>
<gate>
<ID>441</ID>
<type>DE_TO</type>
<position>130,62.5</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-6</lparam></gate>
<gate>
<ID>442</ID>
<type>DE_TO</type>
<position>130,60</position>
<input>
<ID>IN_0</ID>339 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-5</lparam></gate>
<gate>
<ID>443</ID>
<type>DE_TO</type>
<position>130,57.5</position>
<input>
<ID>IN_0</ID>338 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-4</lparam></gate>
<gate>
<ID>444</ID>
<type>DE_TO</type>
<position>130,55</position>
<input>
<ID>IN_0</ID>337 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-3</lparam></gate>
<gate>
<ID>445</ID>
<type>DE_TO</type>
<position>130,52.5</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-2</lparam></gate>
<gate>
<ID>446</ID>
<type>DE_TO</type>
<position>130,50</position>
<input>
<ID>IN_0</ID>335 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-1</lparam></gate>
<gate>
<ID>836</ID>
<type>CC_PULSE</type>
<position>9,30</position>
<output>
<ID>OUT_0</ID>663 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 20</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>455</ID>
<type>AA_LABEL</type>
<position>81,67</position>
<gparam>LABEL_TEXT R0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>456</ID>
<type>AA_LABEL</type>
<position>121.5,67.5</position>
<gparam>LABEL_TEXT R1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>847</ID>
<type>AA_LABEL</type>
<position>40,34</position>
<gparam>LABEL_TEXT Note: issue with timing</gparam>
<gparam>TEXT_HEIGHT 0.1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>462</ID>
<type>DE_TO</type>
<position>-29,43.5</position>
<input>
<ID>IN_0</ID>601 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLOCK-PULSE</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>-15,6</position>
<gparam>LABEL_TEXT Instruction Sequencer</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>465</ID>
<type>DA_FROM</type>
<position>69.5,50</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-1</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>69.5,52.5</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-2</lparam></gate>
<gate>
<ID>467</ID>
<type>DA_FROM</type>
<position>-7.5,48</position>
<input>
<ID>IN_0</ID>354 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID RESET-PC-IN</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>69.5,65</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-7</lparam></gate>
<gate>
<ID>469</ID>
<type>DA_FROM</type>
<position>-17,63</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-PC</lparam></gate>
<gate>
<ID>470</ID>
<type>DA_FROM</type>
<position>69.5,57.5</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-4</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>147,37</position>
<gparam>LABEL_TEXT MBR</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>471</ID>
<type>DA_FROM</type>
<position>-14,65.5</position>
<input>
<ID>IN_0</ID>356 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID INCREMENT-PC</lparam></gate>
<gate>
<ID>472</ID>
<type>DA_FROM</type>
<position>69.5,60</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-5</lparam></gate>
<gate>
<ID>474</ID>
<type>DA_FROM</type>
<position>69.5,62.5</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-6</lparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>113.5,-2</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID REG-SELECT</lparam></gate>
<gate>
<ID>475</ID>
<type>DA_FROM</type>
<position>27,69</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LOAD-IR</lparam></gate>
<gate>
<ID>476</ID>
<type>DA_FROM</type>
<position>69.5,55</position>
<input>
<ID>IN_0</ID>312 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-3</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>-36.5,48.5</position>
<input>
<ID>IN_0</ID>352 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID CLOCK-PULSE-IN</lparam></gate>
<gate>
<ID>477</ID>
<type>DA_FROM</type>
<position>72.5,68</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LOAD-R0</lparam></gate>
<gate>
<ID>478</ID>
<type>DA_FROM</type>
<position>114,68</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LOAD-R1</lparam></gate>
<gate>
<ID>479</ID>
<type>DA_FROM</type>
<position>69.5,47.5</position>
<input>
<ID>IN_0</ID>309 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-0</lparam></gate>
<gate>
<ID>90</ID>
<type>FF_GND</type>
<position>73.5,-1.5</position>
<output>
<ID>OUT_0</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>481</ID>
<type>DA_FROM</type>
<position>111,50</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-1</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>36,2.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LOAD-MAR</lparam></gate>
<gate>
<ID>483</ID>
<type>DA_FROM</type>
<position>111,52.5</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-2</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>89.5,-3.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-2</lparam></gate>
<gate>
<ID>95</ID>
<type>DE_TO</type>
<position>89.5,-6</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-1</lparam></gate>
<gate>
<ID>485</ID>
<type>DA_FROM</type>
<position>111,65</position>
<input>
<ID>IN_0</ID>329 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-7</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>89.5,-8.5</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-0</lparam></gate>
<gate>
<ID>487</ID>
<type>DA_FROM</type>
<position>111,57.5</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-4</lparam></gate>
<gate>
<ID>489</ID>
<type>DA_FROM</type>
<position>111,60</position>
<input>
<ID>IN_0</ID>343 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-5</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>82,5.5</position>
<gparam>LABEL_TEXT OP</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>490</ID>
<type>DA_FROM</type>
<position>45.5,22.5</position>
<input>
<ID>IN_0</ID>368 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-2</lparam></gate>
<gate>
<ID>491</ID>
<type>DA_FROM</type>
<position>45.5,20.5</position>
<input>
<ID>IN_0</ID>366 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-1</lparam></gate>
<gate>
<ID>492</ID>
<type>DA_FROM</type>
<position>45.5,18.5</position>
<input>
<ID>IN_0</ID>367 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-0</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>111,62.5</position>
<input>
<ID>IN_0</ID>330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-6</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_DFF_LOW</type>
<position>108.5,-4</position>
<input>
<ID>IN_0</ID>152 </input>
<output>
<ID>OUT_0</ID>146 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>494</ID>
<type>BE_DECODER_3x8</type>
<position>52,27.5</position>
<input>
<ID>IN_0</ID>367 </input>
<input>
<ID>IN_1</ID>366 </input>
<input>
<ID>IN_2</ID>368 </input>
<output>
<ID>OUT_0</ID>369 </output>
<output>
<ID>OUT_1</ID>370 </output>
<output>
<ID>OUT_2</ID>371 </output>
<output>
<ID>OUT_3</ID>372 </output>
<output>
<ID>OUT_4</ID>373 </output>
<output>
<ID>OUT_5</ID>374 </output>
<output>
<ID>OUT_6</ID>375 </output>
<output>
<ID>OUT_7</ID>376 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_TOGGLE</type>
<position>44,-11</position>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>111,55</position>
<input>
<ID>IN_0</ID>333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-3</lparam></gate>
<gate>
<ID>496</ID>
<type>DA_FROM</type>
<position>111,47.5</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-0</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_TOGGLE</type>
<position>83.5,-12.5</position>
<output>
<ID>OUT_0</ID>163 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>497</ID>
<type>DE_TO</type>
<position>61.5,18</position>
<input>
<ID>IN_0</ID>369 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-STOP</lparam></gate>
<gate>
<ID>498</ID>
<type>DE_TO</type>
<position>61.5,35.5</position>
<input>
<ID>IN_0</ID>376 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-JUMP</lparam></gate>
<gate>
<ID>499</ID>
<type>DE_TO</type>
<position>61.5,33</position>
<input>
<ID>IN_0</ID>375 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-SUB</lparam></gate>
<gate>
<ID>500</ID>
<type>DE_TO</type>
<position>61.5,30.5</position>
<input>
<ID>IN_0</ID>374 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-ADD</lparam></gate>
<gate>
<ID>501</ID>
<type>DE_TO</type>
<position>61.5,28</position>
<input>
<ID>IN_0</ID>373 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-STORE</lparam></gate>
<gate>
<ID>502</ID>
<type>DE_TO</type>
<position>61.5,25.5</position>
<input>
<ID>IN_0</ID>372 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-LOAD</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>79,2</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LOAD-OP</lparam></gate>
<gate>
<ID>503</ID>
<type>DE_TO</type>
<position>61.5,23</position>
<input>
<ID>IN_0</ID>371 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-WRITE</lparam></gate>
<gate>
<ID>504</ID>
<type>DE_TO</type>
<position>61.5,20.5</position>
<input>
<ID>IN_0</ID>370 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-READ</lparam></gate>
<gate>
<ID>115</ID>
<type>DA_FROM</type>
<position>113.5,-11</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID LOAD-REG</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_LABEL</type>
<position>54.5,39.5</position>
<gparam>LABEL_TEXT Instruction Decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_AND2</type>
<position>108.5,-12</position>
<input>
<ID>IN_0</ID>352 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>107,2</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID IR-REG</lparam></gate>
<gate>
<ID>515</ID>
<type>CC_PULSE</type>
<position>-33,43.5</position>
<output>
<ID>OUT_0</ID>601 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>521</ID>
<type>DA_FROM</type>
<position>97,40</position>
<input>
<ID>IN_0</ID>386 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READ-PENDING</lparam></gate>
<gate>
<ID>523</ID>
<type>GA_LED</type>
<position>100.5,40</position>
<input>
<ID>N_in0</ID>386 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>524</ID>
<type>DA_FROM</type>
<position>129.5,40</position>
<input>
<ID>IN_0</ID>387 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OUTPUT-READY</lparam></gate>
<gate>
<ID>525</ID>
<type>GA_LED</type>
<position>132.5,40</position>
<input>
<ID>N_in0</ID>387 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>526</ID>
<type>AA_TOGGLE</type>
<position>81.5,24</position>
<output>
<ID>OUT_0</ID>397 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>527</ID>
<type>AA_TOGGLE</type>
<position>81.5,21.5</position>
<output>
<ID>OUT_0</ID>396 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>528</ID>
<type>AA_TOGGLE</type>
<position>81.5,19</position>
<output>
<ID>OUT_0</ID>395 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>529</ID>
<type>AA_TOGGLE</type>
<position>81.5,16.5</position>
<output>
<ID>OUT_0</ID>394 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>530</ID>
<type>AE_REGISTER8</type>
<position>91.5,24.5</position>
<input>
<ID>IN_0</ID>394 </input>
<input>
<ID>IN_1</ID>395 </input>
<input>
<ID>IN_2</ID>396 </input>
<input>
<ID>IN_3</ID>397 </input>
<input>
<ID>IN_4</ID>398 </input>
<input>
<ID>IN_5</ID>399 </input>
<input>
<ID>IN_6</ID>400 </input>
<input>
<ID>IN_7</ID>401 </input>
<output>
<ID>OUT_0</ID>388 </output>
<output>
<ID>OUT_1</ID>389 </output>
<output>
<ID>OUT_2</ID>403 </output>
<output>
<ID>OUT_3</ID>404 </output>
<output>
<ID>OUT_4</ID>390 </output>
<output>
<ID>OUT_5</ID>391 </output>
<output>
<ID>OUT_6</ID>392 </output>
<output>
<ID>OUT_7</ID>393 </output>
<input>
<ID>clear</ID>362 </input>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>load</ID>402 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>531</ID>
<type>DE_TO</type>
<position>100,16</position>
<input>
<ID>IN_0</ID>388 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-0</lparam></gate>
<gate>
<ID>532</ID>
<type>DE_TO</type>
<position>100,33.5</position>
<input>
<ID>IN_0</ID>393 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-7</lparam></gate>
<gate>
<ID>533</ID>
<type>DE_TO</type>
<position>100,31</position>
<input>
<ID>IN_0</ID>392 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-6</lparam></gate>
<gate>
<ID>534</ID>
<type>DE_TO</type>
<position>100,28.5</position>
<input>
<ID>IN_0</ID>391 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-5</lparam></gate>
<gate>
<ID>535</ID>
<type>DE_TO</type>
<position>100,26</position>
<input>
<ID>IN_0</ID>390 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-4</lparam></gate>
<gate>
<ID>536</ID>
<type>DE_TO</type>
<position>100,23.5</position>
<input>
<ID>IN_0</ID>404 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-3</lparam></gate>
<gate>
<ID>537</ID>
<type>DE_TO</type>
<position>100,21</position>
<input>
<ID>IN_0</ID>403 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-2</lparam></gate>
<gate>
<ID>538</ID>
<type>DE_TO</type>
<position>100,18.5</position>
<input>
<ID>IN_0</ID>389 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-1</lparam></gate>
<gate>
<ID>539</ID>
<type>AA_TOGGLE</type>
<position>81.5,34</position>
<output>
<ID>OUT_0</ID>401 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>540</ID>
<type>AA_TOGGLE</type>
<position>81.5,31.5</position>
<output>
<ID>OUT_0</ID>400 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>541</ID>
<type>AA_TOGGLE</type>
<position>81.5,29</position>
<output>
<ID>OUT_0</ID>399 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>542</ID>
<type>AA_TOGGLE</type>
<position>81.5,26.5</position>
<output>
<ID>OUT_0</ID>398 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>543</ID>
<type>AA_LABEL</type>
<position>94,35.5</position>
<gparam>LABEL_TEXT IN</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>544</ID>
<type>DA_FROM</type>
<position>85,37</position>
<input>
<ID>IN_0</ID>402 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LOAD-IN</lparam></gate>
<gate>
<ID>549</ID>
<type>AA_TOGGLE</type>
<position>-16.5,31.5</position>
<output>
<ID>OUT_0</ID>204 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>550</ID>
<type>AA_TOGGLE</type>
<position>-16.5,29</position>
<output>
<ID>OUT_0</ID>206 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>551</ID>
<type>AA_TOGGLE</type>
<position>-16.5,26.5</position>
<output>
<ID>OUT_0</ID>208 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>556</ID>
<type>AA_TOGGLE</type>
<position>-16.5,24</position>
<output>
<ID>OUT_0</ID>357 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_TOGGLE</type>
<position>-16.5,21.5</position>
<output>
<ID>OUT_0</ID>361 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>564</ID>
<type>AE_REGISTER8</type>
<position>127,24.5</position>
<input>
<ID>IN_0</ID>226 </input>
<input>
<ID>IN_1</ID>229 </input>
<input>
<ID>IN_2</ID>230 </input>
<input>
<ID>IN_3</ID>231 </input>
<input>
<ID>IN_4</ID>232 </input>
<input>
<ID>IN_5</ID>233 </input>
<input>
<ID>IN_6</ID>228 </input>
<input>
<ID>IN_7</ID>227 </input>
<output>
<ID>OUT_0</ID>439 </output>
<output>
<ID>OUT_1</ID>440 </output>
<output>
<ID>OUT_2</ID>441 </output>
<output>
<ID>OUT_3</ID>442 </output>
<output>
<ID>OUT_4</ID>443 </output>
<output>
<ID>OUT_5</ID>444 </output>
<output>
<ID>OUT_6</ID>445 </output>
<output>
<ID>OUT_7</ID>446 </output>
<input>
<ID>clear</ID>363 </input>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>load</ID>438 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>118.5,2</position>
<input>
<ID>N_in2</ID>146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>581</ID>
<type>AA_LABEL</type>
<position>130.5,36.5</position>
<gparam>LABEL_TEXT OUT</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>582</ID>
<type>DA_FROM</type>
<position>120.5,37</position>
<input>
<ID>IN_0</ID>438 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LOAD-OUT</lparam></gate>
<gate>
<ID>584</ID>
<type>GA_LED</type>
<position>135,34</position>
<input>
<ID>N_in0</ID>446 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>585</ID>
<type>GA_LED</type>
<position>135,31.5</position>
<input>
<ID>N_in0</ID>445 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>586</ID>
<type>GA_LED</type>
<position>135,29</position>
<input>
<ID>N_in0</ID>444 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>587</ID>
<type>GA_LED</type>
<position>135,26.5</position>
<input>
<ID>N_in0</ID>443 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>588</ID>
<type>GA_LED</type>
<position>135,24</position>
<input>
<ID>N_in0</ID>442 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>589</ID>
<type>GA_LED</type>
<position>135,21.5</position>
<input>
<ID>N_in0</ID>441 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>590</ID>
<type>GA_LED</type>
<position>135,19</position>
<input>
<ID>N_in0</ID>440 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>591</ID>
<type>GA_LED</type>
<position>135,16.5</position>
<input>
<ID>N_in0</ID>439 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>603</ID>
<type>AA_TOGGLE</type>
<position>-16.5,19</position>
<output>
<ID>OUT_0</ID>377 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>607</ID>
<type>AA_TOGGLE</type>
<position>-16.5,16.5</position>
<output>
<ID>OUT_0</ID>365 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>609</ID>
<type>AA_TOGGLE</type>
<position>-16.5,14</position>
<output>
<ID>OUT_0</ID>364 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>617</ID>
<type>DE_TO</type>
<position>-12.5,31.5</position>
<input>
<ID>IN_0</ID>204 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-REG-USER</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>118,19</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-1</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>118,21.5</position>
<input>
<ID>IN_0</ID>230 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-2</lparam></gate>
<gate>
<ID>230</ID>
<type>DA_FROM</type>
<position>118,34</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-7</lparam></gate>
<gate>
<ID>620</ID>
<type>DE_TO</type>
<position>-12.5,29</position>
<input>
<ID>IN_0</ID>206 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-3-USER</lparam></gate>
<gate>
<ID>231</ID>
<type>DA_FROM</type>
<position>118,26.5</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-4</lparam></gate>
<gate>
<ID>621</ID>
<type>DE_TO</type>
<position>-12.5,26.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-2-USER</lparam></gate>
<gate>
<ID>232</ID>
<type>DA_FROM</type>
<position>118,29</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-5</lparam></gate>
<gate>
<ID>622</ID>
<type>DE_TO</type>
<position>-12.5,24</position>
<input>
<ID>IN_0</ID>357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-1-USER</lparam></gate>
<gate>
<ID>233</ID>
<type>DA_FROM</type>
<position>118,31.5</position>
<input>
<ID>IN_0</ID>228 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-6</lparam></gate>
<gate>
<ID>623</ID>
<type>DE_TO</type>
<position>-12.5,21.5</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-0-USER</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>118,24</position>
<input>
<ID>IN_0</ID>231 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-3</lparam></gate>
<gate>
<ID>624</ID>
<type>DE_TO</type>
<position>-12.5,19</position>
<input>
<ID>IN_0</ID>377 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-2-USER</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>118,16.5</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-0</lparam></gate>
<gate>
<ID>1037</ID>
<type>CC_PULSE</type>
<position>81,43</position>
<output>
<ID>OUT_0</ID>859 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 10</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1039</ID>
<type>DE_TO</type>
<position>85,43</position>
<input>
<ID>IN_0</ID>859 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CONTINUE-PROGRAM</lparam></gate>
<gate>
<ID>276</ID>
<type>DA_FROM</type>
<position>149.5,19</position>
<input>
<ID>IN_0</ID>215 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-1</lparam></gate>
<gate>
<ID>277</ID>
<type>DA_FROM</type>
<position>149.5,21.5</position>
<input>
<ID>IN_0</ID>214 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-2</lparam></gate>
<gate>
<ID>667</ID>
<type>AA_LABEL</type>
<position>24.5,34.5</position>
<gparam>LABEL_TEXT Usage: Must be high to write instruction and low to use instruction ram</gparam>
<gparam>TEXT_HEIGHT 0.6</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>DA_FROM</type>
<position>149.5,24</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-3</lparam></gate>
<gate>
<ID>279</ID>
<type>GA_LED</type>
<position>152.5,34</position>
<input>
<ID>N_in0</ID>209 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>280</ID>
<type>GA_LED</type>
<position>152.5,31.5</position>
<input>
<ID>N_in0</ID>210 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>281</ID>
<type>GA_LED</type>
<position>152.5,29</position>
<input>
<ID>N_in0</ID>211 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>282</ID>
<type>GA_LED</type>
<position>152.5,26.5</position>
<input>
<ID>N_in0</ID>212 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>283</ID>
<type>GA_LED</type>
<position>152.5,24</position>
<input>
<ID>N_in0</ID>213 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>284</ID>
<type>GA_LED</type>
<position>152.5,21.5</position>
<input>
<ID>N_in0</ID>214 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>285</ID>
<type>GA_LED</type>
<position>152.5,19</position>
<input>
<ID>N_in0</ID>215 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>286</ID>
<type>GA_LED</type>
<position>152.5,16.5</position>
<input>
<ID>N_in0</ID>216 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>287</ID>
<type>DA_FROM</type>
<position>149.5,26.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-4</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>149.5,29</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-5</lparam></gate>
<gate>
<ID>289</ID>
<type>DA_FROM</type>
<position>149.5,31.5</position>
<input>
<ID>IN_0</ID>210 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-6</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>149.5,34</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-7</lparam></gate>
<gate>
<ID>291</ID>
<type>DA_FROM</type>
<position>149.5,16.5</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-0</lparam></gate>
<gate>
<ID>1076</ID>
<type>AA_LABEL</type>
<position>-23,39</position>
<gparam>LABEL_TEXT Usage: Press RESET-PC before RUN-PROGRAM</gparam>
<gparam>TEXT_HEIGHT 0.6</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1078</ID>
<type>AA_LABEL</type>
<position>-22,38</position>
<gparam>LABEL_TEXT  to ensure no instructions are missed</gparam>
<gparam>TEXT_HEIGHT 0.6</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>711</ID>
<type>AA_TOGGLE</type>
<position>80.5,48.5</position>
<output>
<ID>OUT_0</ID>553 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>712</ID>
<type>AA_TOGGLE</type>
<position>121.5,48.5</position>
<output>
<ID>OUT_0</ID>554 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>332</ID>
<type>EE_VDD</type>
<position>-19,-5.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>722</ID>
<type>DE_TO</type>
<position>-12.5,16.5</position>
<input>
<ID>IN_0</ID>365 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-1-USER</lparam></gate>
<gate>
<ID>726</ID>
<type>DE_TO</type>
<position>-12.5,14</position>
<input>
<ID>IN_0</ID>364 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-0-USER</lparam></gate>
<gate>
<ID>740</ID>
<type>DA_FROM</type>
<position>25,64</position>
<input>
<ID>IN_0</ID>382 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-REG-IN</lparam></gate>
<gate>
<ID>741</ID>
<type>DA_FROM</type>
<position>25,62</position>
<input>
<ID>IN_0</ID>383 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-3-IN</lparam></gate>
<gate>
<ID>742</ID>
<type>DA_FROM</type>
<position>25,60</position>
<input>
<ID>IN_0</ID>405 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-2-IN</lparam></gate>
<gate>
<ID>743</ID>
<type>DA_FROM</type>
<position>25,58</position>
<input>
<ID>IN_0</ID>515 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-1-IN</lparam></gate>
<gate>
<ID>744</ID>
<type>DA_FROM</type>
<position>25,56</position>
<input>
<ID>IN_0</ID>481 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-0-IN</lparam></gate>
<gate>
<ID>745</ID>
<type>DA_FROM</type>
<position>25,54</position>
<input>
<ID>IN_0</ID>463 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-2-IN</lparam></gate>
<gate>
<ID>746</ID>
<type>DA_FROM</type>
<position>25,52</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-1-IN</lparam></gate>
<gate>
<ID>747</ID>
<type>DA_FROM</type>
<position>25,50</position>
<input>
<ID>IN_0</ID>437 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-0-IN</lparam></gate>
<gate>
<ID>754</ID>
<type>AA_LABEL</type>
<position>9,39.5</position>
<gparam>LABEL_TEXT Instruction Inputs</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>370</ID>
<type>AA_TOGGLE</type>
<position>92.5,18</position>
<output>
<ID>OUT_0</ID>362 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>371</ID>
<type>AA_TOGGLE</type>
<position>128,17.5</position>
<output>
<ID>OUT_0</ID>363 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>386</ID>
<type>AA_REGISTER4</type>
<position>-11,56</position>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>315 </input>
<input>
<ID>IN_2</ID>316 </input>
<input>
<ID>IN_3</ID>317 </input>
<output>
<ID>OUT_0</ID>305 </output>
<output>
<ID>OUT_1</ID>306 </output>
<output>
<ID>OUT_2</ID>307 </output>
<output>
<ID>OUT_3</ID>308 </output>
<input>
<ID>clear</ID>354 </input>
<input>
<ID>clock</ID>352 </input>
<input>
<ID>count_enable</ID>356 </input>
<input>
<ID>count_up</ID>32 </input>
<input>
<ID>load</ID>355 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>387</ID>
<type>AA_LABEL</type>
<position>-7.5,67.5</position>
<gparam>LABEL_TEXT PC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>776</ID>
<type>AA_TOGGLE</type>
<position>9,32.5</position>
<output>
<ID>OUT_0</ID>522 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>386</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>99,40,99.5,40</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<connection>
<GID>523</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,40,131.5,40</points>
<connection>
<GID>524</GID>
<name>IN_0</name></connection>
<connection>
<GID>525</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,16,96,21.5</points>
<intersection>16 4</intersection>
<intersection>21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>95.5,21.5,96,21.5</points>
<connection>
<GID>530</GID>
<name>OUT_0</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>96,16,98,16</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>389</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,18.5,96.5,22.5</points>
<intersection>18.5 1</intersection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,18.5,98,18.5</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,22.5,96.5,22.5</points>
<connection>
<GID>530</GID>
<name>OUT_1</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>390</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,26,98,26</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<intersection>95.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>95.5,25.5,95.5,26</points>
<connection>
<GID>530</GID>
<name>OUT_4</name></connection>
<intersection>26 1</intersection></vsegment></shape></wire>
<wire>
<ID>583</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,-20,-18.5,-17</points>
<connection>
<GID>12</GID>
<name>clear</name></connection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18.5,-20,-17,-20</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>-18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,26.5,97.5,28.5</points>
<intersection>26.5 2</intersection>
<intersection>28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,28.5,98,28.5</points>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,26.5,97.5,26.5</points>
<connection>
<GID>530</GID>
<name>OUT_5</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,27.5,97,31</points>
<intersection>27.5 2</intersection>
<intersection>31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,31,98,31</points>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,27.5,97,27.5</points>
<connection>
<GID>530</GID>
<name>OUT_6</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,28.5,96.5,33.5</points>
<intersection>28.5 2</intersection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,33.5,98,33.5</points>
<connection>
<GID>532</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,28.5,96.5,28.5</points>
<connection>
<GID>530</GID>
<name>OUT_7</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,16.5,87.5,21.5</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>83.5,16.5,87.5,16.5</points>
<connection>
<GID>529</GID>
<name>OUT_0</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,19,86.5,22.5</points>
<intersection>19 2</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,22.5,87.5,22.5</points>
<connection>
<GID>530</GID>
<name>IN_1</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,19,86.5,19</points>
<connection>
<GID>528</GID>
<name>OUT_0</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-3,39,-1</points>
<connection>
<GID>18</GID>
<name>IN_3</name></connection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-1,39,-1</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,21.5,86,23.5</points>
<intersection>21.5 2</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,23.5,87.5,23.5</points>
<connection>
<GID>530</GID>
<name>IN_2</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,21.5,86,21.5</points>
<connection>
<GID>527</GID>
<name>OUT_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,31.5,-14.5,31.5</points>
<connection>
<GID>549</GID>
<name>OUT_0</name></connection>
<connection>
<GID>617</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,24,85.5,24.5</points>
<intersection>24 2</intersection>
<intersection>24.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>83.5,24,85.5,24</points>
<connection>
<GID>526</GID>
<name>OUT_0</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>85.5,24.5,87.5,24.5</points>
<connection>
<GID>530</GID>
<name>IN_3</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-4,38,-3.5</points>
<intersection>-4 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-4,39,-4</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-3.5,38,-3.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,25.5,84.5,26.5</points>
<intersection>25.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,25.5,87.5,25.5</points>
<connection>
<GID>530</GID>
<name>IN_4</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,26.5,84.5,26.5</points>
<connection>
<GID>542</GID>
<name>OUT_0</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-6,38,-5</points>
<intersection>-6 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-5,39,-5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-6,38,-6</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,29,-14.5,29</points>
<connection>
<GID>550</GID>
<name>OUT_0</name></connection>
<connection>
<GID>620</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>399</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,26.5,85,29</points>
<intersection>26.5 1</intersection>
<intersection>29 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,26.5,87.5,26.5</points>
<connection>
<GID>530</GID>
<name>IN_5</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>83.5,29,85,29</points>
<connection>
<GID>541</GID>
<name>OUT_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-8.5,38.5,-6</points>
<intersection>-8.5 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-6,39,-6</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-8.5,38.5,-8.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>400</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,27.5,86,31.5</points>
<intersection>27.5 1</intersection>
<intersection>31.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,27.5,87.5,27.5</points>
<connection>
<GID>530</GID>
<name>IN_6</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>83.5,31.5,86,31.5</points>
<connection>
<GID>540</GID>
<name>OUT_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-3,48,-1</points>
<intersection>-3 2</intersection>
<intersection>-1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-1,49,-1</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-3,48,-3</points>
<connection>
<GID>18</GID>
<name>OUT_3</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-14.5,26.5,-14.5,26.5</points>
<connection>
<GID>551</GID>
<name>OUT_0</name></connection>
<connection>
<GID>621</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>401</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,28.5,87,34</points>
<intersection>28.5 1</intersection>
<intersection>34 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,28.5,87.5,28.5</points>
<connection>
<GID>530</GID>
<name>IN_7</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>83.5,34,87,34</points>
<connection>
<GID>539</GID>
<name>OUT_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-8.5,47.5,-6</points>
<intersection>-8.5 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-6,47.5,-6</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-8.5,49,-8.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,34,151.5,34</points>
<connection>
<GID>279</GID>
<name>N_in0</name></connection>
<connection>
<GID>290</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>402</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,30.5,90.5,37</points>
<connection>
<GID>530</GID>
<name>load</name></connection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,37,90.5,37</points>
<connection>
<GID>544</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-6,48,-5</points>
<intersection>-6 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-5,48,-5</points>
<connection>
<GID>18</GID>
<name>OUT_1</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-6,49,-6</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,31.5,151.5,31.5</points>
<connection>
<GID>280</GID>
<name>N_in0</name></connection>
<connection>
<GID>289</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>403</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,21,97,23.5</points>
<intersection>21 1</intersection>
<intersection>23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,21,98,21</points>
<connection>
<GID>537</GID>
<name>IN_0</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,23.5,97,23.5</points>
<connection>
<GID>530</GID>
<name>OUT_2</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-4,48,-3.5</points>
<intersection>-4 1</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-4,48,-4</points>
<connection>
<GID>18</GID>
<name>OUT_2</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-3.5,49,-3.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,29,151.5,29</points>
<connection>
<GID>281</GID>
<name>N_in0</name></connection>
<connection>
<GID>288</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>404</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,23.5,97.5,24.5</points>
<intersection>23.5 1</intersection>
<intersection>24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97.5,23.5,98,23.5</points>
<connection>
<GID>536</GID>
<name>IN_0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,24.5,97.5,24.5</points>
<connection>
<GID>530</GID>
<name>OUT_3</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,41,-31,41</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>31</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,26.5,151.5,26.5</points>
<connection>
<GID>282</GID>
<name>N_in0</name></connection>
<connection>
<GID>287</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>405</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,58.5,28,60</points>
<intersection>58.5 1</intersection>
<intersection>60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,58.5,29,58.5</points>
<connection>
<GID>392</GID>
<name>IN_5</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,60,28,60</points>
<connection>
<GID>742</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,24,151.5,24</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<connection>
<GID>283</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,21.5,151.5,21.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<connection>
<GID>284</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>-15.5,-11,-14.5,-11</points>
<connection>
<GID>12</GID>
<name>OUT_3</name></connection>
<connection>
<GID>37</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,19,151.5,19</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<connection>
<GID>285</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>601</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,43.5,-31,43.5</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<connection>
<GID>515</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>-15.5,-12,-14.5,-12</points>
<connection>
<GID>12</GID>
<name>OUT_2</name></connection>
<connection>
<GID>37</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151.5,16.5,151.5,16.5</points>
<connection>
<GID>286</GID>
<name>N_in0</name></connection>
<connection>
<GID>291</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>-15.5,-13,-14.5,-13</points>
<connection>
<GID>12</GID>
<name>OUT_1</name></connection>
<connection>
<GID>37</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>6</ID>
<points>-15.5,-14,-14.5,-14</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-17.5,-8,-14</points>
<intersection>-17.5 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-14,-8,-14</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>-8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-17.5,-5,-17.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-15.5,-7.5,-13</points>
<intersection>-15.5 5</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-13,-7.5,-13</points>
<connection>
<GID>37</GID>
<name>OUT_1</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-7.5,-15.5,-5,-15.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-13.5,-7,-12</points>
<intersection>-13.5 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-12,-7,-12</points>
<connection>
<GID>37</GID>
<name>OUT_2</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7,-13.5,-5,-13.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-11.5,-6.5,-11</points>
<intersection>-11.5 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-11,-6.5,-11</points>
<connection>
<GID>37</GID>
<name>OUT_3</name></connection>
<intersection>-6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,-11.5,-5,-11.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-10,-5,-10</points>
<connection>
<GID>37</GID>
<name>OUT_4</name></connection>
<intersection>-5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-5,-10,-5,-9.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-10 1</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-9,-5,-7.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8.5,-9,-5,-9</points>
<connection>
<GID>37</GID>
<name>OUT_5</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-8,-5.5,-5.5</points>
<intersection>-8 2</intersection>
<intersection>-5.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-8,-5.5,-8</points>
<connection>
<GID>37</GID>
<name>OUT_6</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-5.5,-5.5,-5,-5.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-10,62.5,-6.5,62.5</points>
<intersection>-10 4</intersection>
<intersection>-6.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6.5,62.5,-6.5,63.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>62.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-10,61,-10,62.5</points>
<connection>
<GID>386</GID>
<name>count_up</name></connection>
<intersection>62.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,16.5,123,21.5</points>
<connection>
<GID>564</GID>
<name>IN_0</name></connection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>120,16.5,123,16.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-7,-6,-3.5</points>
<intersection>-7 2</intersection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-3.5,-5,-3.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-7,-6,-7</points>
<connection>
<GID>37</GID>
<name>OUT_7</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,28.5,123,34</points>
<connection>
<GID>564</GID>
<name>IN_7</name></connection>
<intersection>34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>120,34,123,34</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-6,-6.5,-1.5</points>
<intersection>-6 2</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,-1.5,-5,-1.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-6,-6.5,-6</points>
<connection>
<GID>37</GID>
<name>OUT_8</name></connection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,27.5,122.5,31.5</points>
<intersection>27.5 1</intersection>
<intersection>31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,27.5,123,27.5</points>
<connection>
<GID>564</GID>
<name>IN_6</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,31.5,122.5,31.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-5,-7,0.5</points>
<intersection>-5 2</intersection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,0.5,-5,0.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-5,-7,-5</points>
<connection>
<GID>37</GID>
<name>OUT_9</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,19,122.5,22.5</points>
<intersection>19 2</intersection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,22.5,123,22.5</points>
<connection>
<GID>564</GID>
<name>IN_1</name></connection>
<intersection>122.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,19,122.5,19</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,21.5,121.5,23.5</points>
<intersection>21.5 2</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,23.5,123,23.5</points>
<connection>
<GID>564</GID>
<name>IN_2</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,21.5,121.5,21.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,24,121.5,24.5</points>
<intersection>24 2</intersection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,24.5,123,24.5</points>
<connection>
<GID>564</GID>
<name>IN_3</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,24,121.5,24</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,25.5,121.5,26.5</points>
<intersection>25.5 1</intersection>
<intersection>26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,25.5,123,25.5</points>
<connection>
<GID>564</GID>
<name>IN_4</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,26.5,121.5,26.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,26.5,122,29</points>
<intersection>26.5 2</intersection>
<intersection>29 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>122,26.5,123,26.5</points>
<connection>
<GID>564</GID>
<name>IN_5</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>120,29,122,29</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire>
<wire>
<ID>627</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,36,-31,36</points>
<connection>
<GID>800</GID>
<name>IN_0</name></connection>
<connection>
<GID>812</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,-8,-19,-6.5</points>
<connection>
<GID>332</GID>
<name>OUT_0</name></connection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,-8,-18.5,-8</points>
<connection>
<GID>12</GID>
<name>count_up</name></connection>
<connection>
<GID>12</GID>
<name>count_enable</name></connection>
<intersection>-19 0</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,50,29,53.5</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>50 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>27,50,29,50</points>
<connection>
<GID>747</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,30.5,126,37</points>
<connection>
<GID>564</GID>
<name>load</name></connection>
<intersection>37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,37,126,37</points>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>439</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,16.5,131,21.5</points>
<connection>
<GID>564</GID>
<name>OUT_0</name></connection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131,16.5,134,16.5</points>
<connection>
<GID>591</GID>
<name>N_in0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>440</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,19,131.5,22.5</points>
<intersection>19 1</intersection>
<intersection>22.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,19,134,19</points>
<connection>
<GID>590</GID>
<name>N_in0</name></connection>
<intersection>131.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,22.5,131.5,22.5</points>
<connection>
<GID>564</GID>
<name>OUT_1</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>441</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,21.5,132,23.5</points>
<intersection>21.5 3</intersection>
<intersection>23.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>131,23.5,132,23.5</points>
<connection>
<GID>564</GID>
<name>OUT_2</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132,21.5,134,21.5</points>
<connection>
<GID>589</GID>
<name>N_in0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>442</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,24,132.5,24.5</points>
<intersection>24 1</intersection>
<intersection>24.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,24,134,24</points>
<connection>
<GID>588</GID>
<name>N_in0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,24.5,132.5,24.5</points>
<connection>
<GID>564</GID>
<name>OUT_3</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>443</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132.5,25.5,132.5,26.5</points>
<intersection>25.5 2</intersection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132.5,26.5,134,26.5</points>
<connection>
<GID>587</GID>
<name>N_in0</name></connection>
<intersection>132.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,25.5,132.5,25.5</points>
<connection>
<GID>564</GID>
<name>OUT_4</name></connection>
<intersection>132.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>444</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>132,26.5,132,29</points>
<intersection>26.5 2</intersection>
<intersection>29 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>131,26.5,132,26.5</points>
<connection>
<GID>564</GID>
<name>OUT_5</name></connection>
<intersection>132 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>132,29,134,29</points>
<connection>
<GID>586</GID>
<name>N_in0</name></connection>
<intersection>132 0</intersection></hsegment></shape></wire>
<wire>
<ID>445</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,27.5,131.5,31.5</points>
<intersection>27.5 3</intersection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>131.5,31.5,134,31.5</points>
<connection>
<GID>585</GID>
<name>N_in0</name></connection>
<intersection>131.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>131,27.5,131.5,27.5</points>
<connection>
<GID>564</GID>
<name>OUT_6</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>446</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,28.5,131,34</points>
<connection>
<GID>564</GID>
<name>OUT_7</name></connection>
<intersection>34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>131,34,134,34</points>
<connection>
<GID>584</GID>
<name>N_in0</name></connection>
<intersection>131 0</intersection></hsegment></shape></wire>
<wire>
<ID>449</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,52,28.5,54.5</points>
<intersection>52 3</intersection>
<intersection>54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,54.5,29,54.5</points>
<connection>
<GID>392</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,52,28.5,52</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,50,115,53.5</points>
<intersection>50 1</intersection>
<intersection>53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,50,115,50</points>
<connection>
<GID>481</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>115,53.5,116.5,53.5</points>
<connection>
<GID>438</GID>
<name>IN_1</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,54,28,55.5</points>
<intersection>54 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,55.5,29,55.5</points>
<connection>
<GID>392</GID>
<name>IN_2</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,54,28,54</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,22,18,22</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,22,18,22</points>
<connection>
<GID>796</GID>
<name>OUT_3</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,16,18,16</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,16,18,16</points>
<connection>
<GID>796</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,20,18,20</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<intersection>20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,20,18,20</points>
<connection>
<GID>796</GID>
<name>OUT_2</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,18,18,18</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,18,18,18</points>
<connection>
<GID>796</GID>
<name>OUT_1</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>663</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,30,11,30</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,30,11,30</points>
<connection>
<GID>836</GID>
<name>OUT_0</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>859</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,43,83,43</points>
<connection>
<GID>1039</GID>
<name>IN_0</name></connection>
<intersection>83 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>83,43,83,43</points>
<connection>
<GID>1037</GID>
<name>OUT_0</name></connection>
<intersection>43 0</intersection></vsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,47.5,116.5,52.5</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>113,47.5,116.5,47.5</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,48,37.5,53.5</points>
<intersection>48 1</intersection>
<intersection>53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,48,39.5,48</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,53.5,37.5,53.5</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,50.5,38,54.5</points>
<intersection>50.5 1</intersection>
<intersection>54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,50.5,39.5,50.5</points>
<connection>
<GID>401</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,54.5,38,54.5</points>
<connection>
<GID>392</GID>
<name>OUT_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>481</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,56,28,56.5</points>
<intersection>56 2</intersection>
<intersection>56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,56.5,29,56.5</points>
<connection>
<GID>392</GID>
<name>IN_3</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,56,28,56</points>
<connection>
<GID>744</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,58,39.5,58</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>37 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>37,57.5,37,58</points>
<connection>
<GID>392</GID>
<name>OUT_4</name></connection>
<intersection>58 1</intersection></vsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,58.5,39,60.5</points>
<intersection>58.5 2</intersection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,60.5,39.5,60.5</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,58.5,39,58.5</points>
<connection>
<GID>392</GID>
<name>OUT_5</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,59.5,38.5,63</points>
<intersection>59.5 2</intersection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,63,39.5,63</points>
<connection>
<GID>396</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,59.5,38.5,59.5</points>
<connection>
<GID>392</GID>
<name>OUT_6</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,60.5,38,65.5</points>
<intersection>60.5 2</intersection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,65.5,39.5,65.5</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,60.5,38,60.5</points>
<connection>
<GID>392</GID>
<name>OUT_7</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,59.5,75.5,65</points>
<connection>
<GID>421</GID>
<name>IN_7</name></connection>
<intersection>65 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>71.5,65,75.5,65</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,52.5,-6,55</points>
<intersection>52.5 1</intersection>
<intersection>55 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,52.5,-5,52.5</points>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-7,55,-6,55</points>
<connection>
<GID>386</GID>
<name>OUT_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,55,-5.5,56</points>
<intersection>55 3</intersection>
<intersection>56 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7,56,-5.5,56</points>
<connection>
<GID>386</GID>
<name>OUT_1</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-5.5,55,-5,55</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,57,-6,57.5</points>
<intersection>57 3</intersection>
<intersection>57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,57.5,-5,57.5</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-7,57,-6,57</points>
<connection>
<GID>386</GID>
<name>OUT_2</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,58,-6,60</points>
<intersection>58 3</intersection>
<intersection>60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,60,-5,60</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-7,58,-6,58</points>
<connection>
<GID>386</GID>
<name>OUT_3</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,47.5,75.5,52.5</points>
<connection>
<GID>421</GID>
<name>IN_0</name></connection>
<intersection>47.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>71.5,47.5,75.5,47.5</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,50,74.5,53.5</points>
<intersection>50 2</intersection>
<intersection>53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,53.5,75.5,53.5</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,50,74.5,50</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,52.5,73.5,54.5</points>
<intersection>52.5 3</intersection>
<intersection>54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,54.5,75.5,54.5</points>
<connection>
<GID>421</GID>
<name>IN_2</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>71.5,52.5,73.5,52.5</points>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,55,73.5,55.5</points>
<intersection>55 3</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,55.5,75.5,55.5</points>
<connection>
<GID>421</GID>
<name>IN_3</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>71.5,55,73.5,55</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,56.5,73.5,57.5</points>
<intersection>56.5 1</intersection>
<intersection>57.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,56.5,75.5,56.5</points>
<connection>
<GID>421</GID>
<name>IN_4</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>71.5,57.5,73.5,57.5</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,52.5,-15,55</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,52.5,-15,52.5</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15.5,55,-15.5,56</points>
<intersection>55 3</intersection>
<intersection>56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15.5,56,-15,56</points>
<connection>
<GID>386</GID>
<name>IN_1</name></connection>
<intersection>-15.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16,55,-15.5,55</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>-15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16,57.5,-15,57.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>-15 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-15,57,-15,57.5</points>
<connection>
<GID>386</GID>
<name>IN_2</name></connection>
<intersection>57.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-15,58,-15,60</points>
<connection>
<GID>386</GID>
<name>IN_3</name></connection>
<intersection>60 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-16,60,-15,60</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<intersection>-15 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,47.5,84,52.5</points>
<intersection>47.5 1</intersection>
<intersection>52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,47.5,87,47.5</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,52.5,84,52.5</points>
<connection>
<GID>421</GID>
<name>OUT_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,50,85,53.5</points>
<intersection>50 1</intersection>
<intersection>53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,50,87,50</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,53.5,85,53.5</points>
<connection>
<GID>421</GID>
<name>OUT_1</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,52.5,85.5,54.5</points>
<intersection>52.5 1</intersection>
<intersection>54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,52.5,87,52.5</points>
<connection>
<GID>428</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,54.5,85.5,54.5</points>
<connection>
<GID>421</GID>
<name>OUT_2</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,55,85,55.5</points>
<intersection>55 1</intersection>
<intersection>55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,55,87,55</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,55.5,85,55.5</points>
<connection>
<GID>421</GID>
<name>OUT_3</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,56.5,86.5,57.5</points>
<intersection>56.5 2</intersection>
<intersection>57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,57.5,87,57.5</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,56.5,86.5,56.5</points>
<connection>
<GID>421</GID>
<name>OUT_4</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>515</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,57.5,28,58</points>
<intersection>57.5 1</intersection>
<intersection>58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,57.5,29,57.5</points>
<connection>
<GID>392</GID>
<name>IN_4</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,58,28,58</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,57.5,86,60</points>
<intersection>57.5 2</intersection>
<intersection>60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,60,87,60</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,57.5,86,57.5</points>
<connection>
<GID>421</GID>
<name>OUT_5</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,58.5,85,62.5</points>
<intersection>58.5 2</intersection>
<intersection>62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,62.5,87,62.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,58.5,85,58.5</points>
<connection>
<GID>421</GID>
<name>OUT_6</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,59.5,84,65</points>
<intersection>59.5 2</intersection>
<intersection>65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,65,87,65</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83.5,59.5,84,59.5</points>
<connection>
<GID>421</GID>
<name>OUT_7</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,57.5,74,60</points>
<intersection>57.5 1</intersection>
<intersection>60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,57.5,75.5,57.5</points>
<connection>
<GID>421</GID>
<name>IN_5</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,60,74,60</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,58.5,74.5,62.5</points>
<intersection>58.5 1</intersection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,58.5,75.5,58.5</points>
<connection>
<GID>421</GID>
<name>IN_6</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,62.5,74.5,62.5</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,59.5,116.5,65</points>
<connection>
<GID>438</GID>
<name>IN_7</name></connection>
<intersection>65 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>113,65,116.5,65</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>522</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>11,32.5,11,32.5</points>
<connection>
<GID>780</GID>
<name>IN_0</name></connection>
<connection>
<GID>776</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,58.5,115.5,62.5</points>
<intersection>58.5 1</intersection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,58.5,116.5,58.5</points>
<connection>
<GID>438</GID>
<name>IN_6</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113,62.5,115.5,62.5</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-8,78,-7</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-7,78.5,-7</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-6,78.5,-6</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>332</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,52.5,114.5,54.5</points>
<intersection>52.5 3</intersection>
<intersection>54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,54.5,116.5,54.5</points>
<connection>
<GID>438</GID>
<name>IN_2</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>113,52.5,114.5,52.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-5,78,-4</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-5,78.5,-5</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,55,114.5,55.5</points>
<intersection>55 3</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,55.5,116.5,55.5</points>
<connection>
<GID>438</GID>
<name>IN_3</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>113,55,114.5,55</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-4,78.5,-0.5</points>
<connection>
<GID>29</GID>
<name>IN_3</name></connection>
<intersection>-0.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-0.5,78.5,-0.5</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,47.5,125,52.5</points>
<intersection>47.5 1</intersection>
<intersection>52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,47.5,128,47.5</points>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,52.5,125,52.5</points>
<connection>
<GID>438</GID>
<name>OUT_0</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,0,42,2.5</points>
<connection>
<GID>18</GID>
<name>load</name></connection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,2.5,42,2.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,50,126,53.5</points>
<intersection>50 1</intersection>
<intersection>53.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,50,128,50</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,53.5,126,53.5</points>
<connection>
<GID>438</GID>
<name>OUT_1</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,52.5,126.5,54.5</points>
<intersection>52.5 1</intersection>
<intersection>54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126.5,52.5,128,52.5</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>126.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,54.5,126.5,54.5</points>
<connection>
<GID>438</GID>
<name>OUT_2</name></connection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-8.5,87,-7</points>
<intersection>-8.5 3</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-7,87,-7</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>87,-8.5,87.5,-8.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,55,126,55.5</points>
<intersection>55 1</intersection>
<intersection>55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,55,128,55</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,55.5,126,55.5</points>
<connection>
<GID>438</GID>
<name>OUT_3</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>86.5,-6,87.5,-6</points>
<connection>
<GID>29</GID>
<name>OUT_1</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,56.5,127.5,57.5</points>
<intersection>56.5 2</intersection>
<intersection>57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,57.5,128,57.5</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,56.5,127.5,56.5</points>
<connection>
<GID>438</GID>
<name>OUT_4</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-5,87,-3.5</points>
<intersection>-5 2</intersection>
<intersection>-3.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>86.5,-5,87,-5</points>
<connection>
<GID>29</GID>
<name>OUT_2</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>87,-3.5,87.5,-3.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-2,112,0</points>
<intersection>-2 3</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112,0,118.5,0</points>
<intersection>112 0</intersection>
<intersection>118.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>111.5,-2,112,-2</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>118.5,0,118.5,1</points>
<connection>
<GID>184</GID>
<name>N_in2</name></connection>
<intersection>0 2</intersection></vsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,57.5,127,60</points>
<intersection>57.5 2</intersection>
<intersection>60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,60,128,60</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,57.5,127,57.5</points>
<connection>
<GID>438</GID>
<name>OUT_5</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,58.5,126,62.5</points>
<intersection>58.5 2</intersection>
<intersection>62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,62.5,128,62.5</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,58.5,126,58.5</points>
<connection>
<GID>438</GID>
<name>OUT_6</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>341</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,59.5,125,65</points>
<intersection>59.5 2</intersection>
<intersection>65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,65,128,65</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,59.5,125,59.5</points>
<connection>
<GID>438</GID>
<name>OUT_7</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-12,105.5,-5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<connection>
<GID>104</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>342</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,56.5,114.5,57.5</points>
<intersection>56.5 1</intersection>
<intersection>57.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,56.5,116.5,56.5</points>
<connection>
<GID>438</GID>
<name>IN_4</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>113,57.5,114.5,57.5</points>
<connection>
<GID>487</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>343</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,57.5,115,60</points>
<intersection>57.5 1</intersection>
<intersection>60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,57.5,116.5,57.5</points>
<connection>
<GID>438</GID>
<name>IN_5</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113,60,115,60</points>
<connection>
<GID>489</GID>
<name>IN_0</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-1,81.5,2</points>
<connection>
<GID>29</GID>
<name>load</name></connection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,2,81.5,2</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-11,111.5,-11</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>118</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-2,105,2</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-2,105.5,-2</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>44,-9,44,-9</points>
<connection>
<GID>18</GID>
<name>clear</name></connection>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>352</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,45.5,-12,52</points>
<connection>
<GID>386</GID>
<name>clock</name></connection>
<intersection>45.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-36.5,45.5,119.5,45.5</points>
<intersection>-36.5 9</intersection>
<intersection>-12 0</intersection>
<intersection>32 4</intersection>
<intersection>78.5 6</intersection>
<intersection>119.5 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>32,45.5,32,51.5</points>
<connection>
<GID>392</GID>
<name>clock</name></connection>
<intersection>45.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>78.5,45.5,78.5,50.5</points>
<connection>
<GID>421</GID>
<name>clock</name></connection>
<intersection>45.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>119.5,45.5,119.5,50.5</points>
<connection>
<GID>438</GID>
<name>clock</name></connection>
<intersection>45.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-36.5,-23.5,-36.5,46.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-23.5 20</intersection>
<intersection>8 10</intersection>
<intersection>45.5 2</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-36.5,8,126,8</points>
<intersection>-36.5 9</intersection>
<intersection>90.5 11</intersection>
<intersection>126 15</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>90.5,8,90.5,19.5</points>
<connection>
<GID>530</GID>
<name>clock</name></connection>
<intersection>8 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>126,8,126,19.5</points>
<connection>
<GID>564</GID>
<name>clock</name></connection>
<intersection>8 10</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-36.5,-23.5,114,-23.5</points>
<intersection>-36.5 9</intersection>
<intersection>-20.5 48</intersection>
<intersection>42 23</intersection>
<intersection>81.5 22</intersection>
<intersection>114 28</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>81.5,-23.5,81.5,-10</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<intersection>-23.5 20</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>42,-23.5,42,-9</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<intersection>-23.5 20</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>114,-23.5,114,-13</points>
<intersection>-23.5 20</intersection>
<intersection>-13 29</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>111.5,-13,114,-13</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>114 28</intersection></hsegment>
<vsegment>
<ID>48</ID>
<points>-20.5,-23.5,-20.5,-17</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>-23.5 20</intersection></vsegment></shape></wire>
<wire>
<ID>354</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,48,-10,52</points>
<connection>
<GID>386</GID>
<name>clear</name></connection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-10,48,-9.5,48</points>
<connection>
<GID>467</GID>
<name>IN_0</name></connection>
<intersection>-10 0</intersection></hsegment></shape></wire>
<wire>
<ID>355</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,61,-12,63</points>
<connection>
<GID>386</GID>
<name>load</name></connection>
<intersection>63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,63,-12,63</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>356</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,61,-11,65.5</points>
<connection>
<GID>386</GID>
<name>count_enable</name></connection>
<intersection>65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,65.5,-11,65.5</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-10.5,83.5,-10</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<connection>
<GID>29</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>357</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,24,-14.5,24</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,24,-14.5,24</points>
<connection>
<GID>556</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,62.5,32,69</points>
<connection>
<GID>392</GID>
<name>load</name></connection>
<intersection>69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,69,32,69</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,61.5,77,68</points>
<intersection>61.5 2</intersection>
<intersection>68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,68,77,68</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,61.5,78.5,61.5</points>
<connection>
<GID>421</GID>
<name>load</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,61.5,118,68</points>
<intersection>61.5 2</intersection>
<intersection>68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,68,118,68</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>118,61.5,119.5,61.5</points>
<connection>
<GID>438</GID>
<name>load</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>553</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>80.5,50.5,80.5,50.5</points>
<connection>
<GID>421</GID>
<name>clear</name></connection>
<connection>
<GID>711</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,21.5,-14.5,21.5</points>
<connection>
<GID>558</GID>
<name>OUT_0</name></connection>
<connection>
<GID>623</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>554</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,50.5,121.5,50.5</points>
<connection>
<GID>438</GID>
<name>clear</name></connection>
<connection>
<GID>712</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>8</ID>
<points>92.5,19.5,92.5,20</points>
<connection>
<GID>370</GID>
<name>OUT_0</name></connection>
<connection>
<GID>530</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>128,19.5,128,19.5</points>
<connection>
<GID>564</GID>
<name>clear</name></connection>
<connection>
<GID>371</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,14,-14.5,14</points>
<connection>
<GID>726</GID>
<name>IN_0</name></connection>
<intersection>14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14.5,14,-14.5,14</points>
<connection>
<GID>609</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-14.5,16.5,-14.5,16.5</points>
<connection>
<GID>607</GID>
<name>OUT_0</name></connection>
<connection>
<GID>722</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,20.5,48.5,20.5</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<intersection>48.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>48.5,20.5,48.5,25</points>
<intersection>20.5 1</intersection>
<intersection>25 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>48.5,25,49,25</points>
<connection>
<GID>494</GID>
<name>IN_1</name></connection>
<intersection>48.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,18.5,49,24</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>18.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,18.5,49,18.5</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,22.5,48,26</points>
<intersection>22.5 6</intersection>
<intersection>26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,26,49,26</points>
<connection>
<GID>494</GID>
<name>IN_2</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>47.5,22.5,48,22.5</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,18,55,24</points>
<connection>
<GID>494</GID>
<name>OUT_0</name></connection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,18,59.5,18</points>
<connection>
<GID>497</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,20.5,56,25</points>
<intersection>20.5 1</intersection>
<intersection>25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,20.5,59.5,20.5</points>
<connection>
<GID>504</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,25,56,25</points>
<connection>
<GID>494</GID>
<name>OUT_1</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,23,57,26</points>
<intersection>23 3</intersection>
<intersection>26 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,26,57,26</points>
<connection>
<GID>494</GID>
<name>OUT_2</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>57,23,59.5,23</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,25.5,57.5,27</points>
<intersection>25.5 4</intersection>
<intersection>27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,27,57.5,27</points>
<connection>
<GID>494</GID>
<name>OUT_3</name></connection>
<intersection>57.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>57.5,25.5,59.5,25.5</points>
<connection>
<GID>502</GID>
<name>IN_0</name></connection>
<intersection>57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,28,59.5,28</points>
<connection>
<GID>494</GID>
<name>OUT_4</name></connection>
<connection>
<GID>501</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>374</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,29,57,30.5</points>
<intersection>29 2</intersection>
<intersection>30.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,29,57,29</points>
<connection>
<GID>494</GID>
<name>OUT_5</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>57,30.5,59.5,30.5</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,30,56.5,33</points>
<intersection>30 2</intersection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,33,59.5,33</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,30,56.5,30</points>
<connection>
<GID>494</GID>
<name>OUT_6</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>376</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,31,55.5,35.5</points>
<intersection>31 2</intersection>
<intersection>35.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,31,55.5,31</points>
<connection>
<GID>494</GID>
<name>OUT_7</name></connection>
<intersection>55.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>55.5,35.5,59.5,35.5</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>377</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14.5,19,-14.5,19</points>
<connection>
<GID>603</GID>
<name>OUT_0</name></connection>
<connection>
<GID>624</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>382</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,60.5,29,64</points>
<connection>
<GID>392</GID>
<name>IN_7</name></connection>
<intersection>64 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>27,64,29,64</points>
<connection>
<GID>740</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>383</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,59.5,28.5,62</points>
<intersection>59.5 1</intersection>
<intersection>62 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,59.5,29,59.5</points>
<connection>
<GID>392</GID>
<name>IN_6</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>27,62,28.5,62</points>
<connection>
<GID>741</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>384</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,53,38.5,55.5</points>
<intersection>53 1</intersection>
<intersection>55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,53,39.5,53</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,55.5,38.5,55.5</points>
<connection>
<GID>392</GID>
<name>OUT_2</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>385</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,55.5,39,56.5</points>
<intersection>55.5 1</intersection>
<intersection>56.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,55.5,39.5,55.5</points>
<connection>
<GID>399</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,56.5,39,56.5</points>
<connection>
<GID>392</GID>
<name>OUT_3</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-305.529,75.6242,-89.6239,-33.5131</PageViewport>
<gate>
<ID>389</ID>
<type>AA_MUX_2x1</type>
<position>-227.5,-44.5</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>625 </input>
<output>
<ID>OUT</ID>118 </output>
<input>
<ID>SEL_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>-194,8</position>
<input>
<ID>IN_0</ID>530 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID WRITE-INSTRUCTION</lparam></gate>
<gate>
<ID>241</ID>
<type>DE_TO</type>
<position>-185,-45.5</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-0-IN</lparam></gate>
<gate>
<ID>629</ID>
<type>AA_MUX_2x1</type>
<position>-225,27</position>
<input>
<ID>IN_0</ID>568 </input>
<input>
<ID>IN_1</ID>435 </input>
<output>
<ID>OUT</ID>426 </output>
<input>
<ID>SEL_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>630</ID>
<type>VA_NMOS</type>
<position>-206,65</position>
<input>
<ID>T_ctrl</ID>434 </input>
<input>
<ID>T_in</ID>549 </input>
<input>
<ID>T_in2</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>632</ID>
<type>VA_NMOS</type>
<position>-203,65</position>
<input>
<ID>T_ctrl</ID>434 </input>
<input>
<ID>T_in</ID>550 </input>
<input>
<ID>T_in2</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>633</ID>
<type>VA_NMOS</type>
<position>-200,65</position>
<input>
<ID>T_ctrl</ID>434 </input>
<input>
<ID>T_in</ID>551 </input>
<input>
<ID>T_in2</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>826</ID>
<type>DA_FROM</type>
<position>-241.5,-13.5</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-REG-USER</lparam></gate>
<gate>
<ID>634</ID>
<type>VA_NMOS</type>
<position>-197,65</position>
<input>
<ID>T_ctrl</ID>434 </input>
<input>
<ID>T_in</ID>552 </input>
<input>
<ID>T_in2</ID>545 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>827</ID>
<type>DA_FROM</type>
<position>-241,-18.5</position>
<input>
<ID>IN_0</ID>619 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-3-USER</lparam></gate>
<gate>
<ID>635</ID>
<type>VA_NMOS</type>
<position>-194,65</position>
<input>
<ID>T_ctrl</ID>434 </input>
<input>
<ID>T_in</ID>557 </input>
<input>
<ID>T_in2</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>636</ID>
<type>VA_NMOS</type>
<position>-191,65</position>
<input>
<ID>T_ctrl</ID>434 </input>
<input>
<ID>T_in</ID>560 </input>
<input>
<ID>T_in2</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>829</ID>
<type>DA_FROM</type>
<position>-241,-23.5</position>
<input>
<ID>IN_0</ID>620 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-2-USER</lparam></gate>
<gate>
<ID>830</ID>
<type>DA_FROM</type>
<position>-241,-28.5</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-1-USER</lparam></gate>
<gate>
<ID>638</ID>
<type>VA_NMOS</type>
<position>-188,65</position>
<input>
<ID>T_ctrl</ID>434 </input>
<input>
<ID>T_in</ID>568 </input>
<input>
<ID>T_in2</ID>578 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>832</ID>
<type>DA_FROM</type>
<position>-241,-33.5</position>
<input>
<ID>IN_0</ID>622 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-0-USER</lparam></gate>
<gate>
<ID>833</ID>
<type>DA_FROM</type>
<position>-241,-38.5</position>
<input>
<ID>IN_0</ID>623 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-2-USER</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_MUX_2x1</type>
<position>-227.5,-49.5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>624 </input>
<output>
<ID>OUT</ID>199 </output>
<input>
<ID>SEL_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>834</ID>
<type>DA_FROM</type>
<position>-241,-43.5</position>
<input>
<ID>IN_0</ID>625 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-1-USER</lparam></gate>
<gate>
<ID>835</ID>
<type>DA_FROM</type>
<position>-241,-48.5</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-0-USER</lparam></gate>
<gate>
<ID>65</ID>
<type>VA_NMOS</type>
<position>-208.5,-11.5</position>
<input>
<ID>T_ctrl</ID>109 </input>
<input>
<ID>T_in</ID>120 </input>
<input>
<ID>T_in2</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>453</ID>
<type>DA_FROM</type>
<position>-238,48</position>
<input>
<ID>IN_0</ID>430 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-IN-4</lparam></gate>
<gate>
<ID>67</ID>
<type>VA_NMOS</type>
<position>-205.5,-11.5</position>
<input>
<ID>T_ctrl</ID>109 </input>
<input>
<ID>T_in</ID>121 </input>
<input>
<ID>T_in2</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>-238,53</position>
<input>
<ID>IN_0</ID>428 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-IN-5</lparam></gate>
<gate>
<ID>69</ID>
<type>VA_NMOS</type>
<position>-202.5,-11.5</position>
<input>
<ID>T_ctrl</ID>109 </input>
<input>
<ID>T_in</ID>123 </input>
<input>
<ID>T_in2</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>-178.5,-14</position>
<gparam>LABEL_TEXT Output Instruction</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>70</ID>
<type>VA_NMOS</type>
<position>-199.5,-11.5</position>
<input>
<ID>T_ctrl</ID>109 </input>
<input>
<ID>T_in</ID>124 </input>
<input>
<ID>T_in2</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>-238,58</position>
<input>
<ID>IN_0</ID>427 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-IN-6</lparam></gate>
<gate>
<ID>71</ID>
<type>VA_NMOS</type>
<position>-196.5,-11.5</position>
<input>
<ID>T_ctrl</ID>109 </input>
<input>
<ID>T_in</ID>125 </input>
<input>
<ID>T_in2</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>458</ID>
<type>DA_FROM</type>
<position>-238,63</position>
<input>
<ID>IN_0</ID>417 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-IN-7</lparam></gate>
<gate>
<ID>460</ID>
<type>AE_REGISTER8</type>
<position>-211,45</position>
<input>
<ID>IN_0</ID>426 </input>
<input>
<ID>IN_1</ID>425 </input>
<input>
<ID>IN_2</ID>424 </input>
<input>
<ID>IN_3</ID>423 </input>
<input>
<ID>IN_4</ID>422 </input>
<input>
<ID>IN_5</ID>421 </input>
<input>
<ID>IN_6</ID>419 </input>
<input>
<ID>IN_7</ID>418 </input>
<output>
<ID>OUT_0</ID>578 </output>
<output>
<ID>OUT_1</ID>547 </output>
<output>
<ID>OUT_2</ID>546 </output>
<output>
<ID>OUT_3</ID>545 </output>
<output>
<ID>OUT_4</ID>544 </output>
<output>
<ID>OUT_5</ID>543 </output>
<output>
<ID>OUT_6</ID>542 </output>
<output>
<ID>OUT_7</ID>436 </output>
<input>
<ID>clear</ID>579 </input>
<input>
<ID>clock</ID>572 </input>
<input>
<ID>load</ID>2 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>461</ID>
<type>DA_FROM</type>
<position>-188,79.5</position>
<input>
<ID>IN_0</ID>434 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID RAM-WRITE</lparam></gate>
<gate>
<ID>75</ID>
<type>VA_NMOS</type>
<position>-193.5,-11.5</position>
<input>
<ID>T_ctrl</ID>109 </input>
<input>
<ID>T_in</ID>129 </input>
<input>
<ID>T_in2</ID>118 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>76</ID>
<type>VA_NMOS</type>
<position>-190.5,-11.5</position>
<input>
<ID>T_ctrl</ID>109 </input>
<input>
<ID>T_in</ID>132 </input>
<input>
<ID>T_in2</ID>199 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>464</ID>
<type>VA_NMOS</type>
<position>-209,65</position>
<input>
<ID>T_ctrl</ID>434 </input>
<input>
<ID>T_in</ID>548 </input>
<input>
<ID>T_in2</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>473</ID>
<type>AA_MUX_2x1</type>
<position>-225,62</position>
<input>
<ID>IN_0</ID>548 </input>
<input>
<ID>IN_1</ID>417 </input>
<output>
<ID>OUT</ID>418 </output>
<input>
<ID>SEL_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>482</ID>
<type>FF_GND</type>
<position>-232.5,88</position>
<output>
<ID>OUT_0</ID>573 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>484</ID>
<type>DA_FROM</type>
<position>-235.5,82.5</position>
<input>
<ID>IN_0</ID>569 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-2</lparam></gate>
<gate>
<ID>98</ID>
<type>VA_NMOS</type>
<position>-211.5,-11.5</position>
<input>
<ID>T_ctrl</ID>109 </input>
<input>
<ID>T_in</ID>119 </input>
<input>
<ID>T_in2</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam></gate>
<gate>
<ID>678</ID>
<type>DA_FROM</type>
<position>-207,87</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CLOCK-PULSE-IN</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_MUX_2x1</type>
<position>-227.5,-14.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>618 </input>
<output>
<ID>OUT</ID>112 </output>
<input>
<ID>SEL_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>486</ID>
<type>EE_VDD</type>
<position>-200,80.5</position>
<output>
<ID>OUT_0</ID>577 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>679</ID>
<type>AE_RAM_8x8</type>
<position>-217,81</position>
<input>
<ID>ADDRESS_0</ID>420 </input>
<input>
<ID>ADDRESS_1</ID>558 </input>
<input>
<ID>ADDRESS_2</ID>569 </input>
<input>
<ID>ADDRESS_3</ID>570 </input>
<input>
<ID>ADDRESS_4</ID>573 </input>
<input>
<ID>ADDRESS_5</ID>573 </input>
<input>
<ID>ADDRESS_6</ID>573 </input>
<input>
<ID>ADDRESS_7</ID>573 </input>
<input>
<ID>DATA_IN_0</ID>568 </input>
<input>
<ID>DATA_IN_1</ID>560 </input>
<input>
<ID>DATA_IN_2</ID>557 </input>
<input>
<ID>DATA_IN_3</ID>552 </input>
<input>
<ID>DATA_IN_4</ID>551 </input>
<input>
<ID>DATA_IN_5</ID>550 </input>
<input>
<ID>DATA_IN_6</ID>549 </input>
<input>
<ID>DATA_IN_7</ID>548 </input>
<output>
<ID>DATA_OUT_0</ID>568 </output>
<output>
<ID>DATA_OUT_1</ID>560 </output>
<output>
<ID>DATA_OUT_2</ID>557 </output>
<output>
<ID>DATA_OUT_3</ID>552 </output>
<output>
<ID>DATA_OUT_4</ID>551 </output>
<output>
<ID>DATA_OUT_5</ID>550 </output>
<output>
<ID>DATA_OUT_6</ID>549 </output>
<output>
<ID>DATA_OUT_7</ID>548 </output>
<input>
<ID>ENABLE_0</ID>577 </input>
<input>
<ID>write_clock</ID>572 </input>
<input>
<ID>write_enable</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 3</lparam>
<lparam>Address:1 2</lparam>
<lparam>Address:12 86</lparam>
<lparam>Address:13 4</lparam>
<lparam>Address:14 2</lparam>
<lparam>Address:15 2</lparam></gate>
<gate>
<ID>680</ID>
<type>AA_LABEL</type>
<position>-214.5,93</position>
<gparam>LABEL_TEXT 16 x 8-bit RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>FF_GND</type>
<position>-235,11.5</position>
<output>
<ID>OUT_0</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>488</ID>
<type>DA_FROM</type>
<position>-238,28</position>
<input>
<ID>IN_0</ID>435 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-IN-0</lparam></gate>
<gate>
<ID>681</ID>
<type>DE_TO</type>
<position>-182.5,59</position>
<input>
<ID>IN_0</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-7</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>-238,6</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-RAM-2</lparam></gate>
<gate>
<ID>682</ID>
<type>DE_TO</type>
<position>-182.5,55</position>
<input>
<ID>IN_0</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-6</lparam></gate>
<gate>
<ID>683</ID>
<type>DE_TO</type>
<position>-182.5,51</position>
<input>
<ID>IN_0</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-5</lparam></gate>
<gate>
<ID>684</ID>
<type>DE_TO</type>
<position>-182.5,47</position>
<input>
<ID>IN_0</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-4</lparam></gate>
<gate>
<ID>685</ID>
<type>DE_TO</type>
<position>-182.5,43</position>
<input>
<ID>IN_0</ID>545 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-3</lparam></gate>
<gate>
<ID>686</ID>
<type>DE_TO</type>
<position>-182.5,39</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-2</lparam></gate>
<gate>
<ID>687</ID>
<type>DE_TO</type>
<position>-182.5,35</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-1</lparam></gate>
<gate>
<ID>688</ID>
<type>DE_TO</type>
<position>-182.5,31</position>
<input>
<ID>IN_0</ID>578 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-0</lparam></gate>
<gate>
<ID>689</ID>
<type>AA_LABEL</type>
<position>-176,62.5</position>
<gparam>LABEL_TEXT Output Bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>110</ID>
<type>DA_FROM</type>
<position>-202,10.5</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CLOCK-PULSE-IN</lparam></gate>
<gate>
<ID>690</ID>
<type>AA_LABEL</type>
<position>-242.5,66</position>
<gparam>LABEL_TEXT Input Bus</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>111</ID>
<type>AE_RAM_8x8</type>
<position>-219.5,4.5</position>
<input>
<ID>ADDRESS_0</ID>669 </input>
<input>
<ID>ADDRESS_1</ID>128 </input>
<input>
<ID>ADDRESS_2</ID>136 </input>
<input>
<ID>ADDRESS_3</ID>148 </input>
<input>
<ID>ADDRESS_4</ID>195 </input>
<input>
<ID>ADDRESS_5</ID>195 </input>
<input>
<ID>ADDRESS_6</ID>195 </input>
<input>
<ID>ADDRESS_7</ID>195 </input>
<input>
<ID>DATA_IN_0</ID>132 </input>
<input>
<ID>DATA_IN_1</ID>129 </input>
<input>
<ID>DATA_IN_2</ID>125 </input>
<input>
<ID>DATA_IN_3</ID>124 </input>
<input>
<ID>DATA_IN_4</ID>123 </input>
<input>
<ID>DATA_IN_5</ID>121 </input>
<input>
<ID>DATA_IN_6</ID>120 </input>
<input>
<ID>DATA_IN_7</ID>119 </input>
<output>
<ID>DATA_OUT_0</ID>132 </output>
<output>
<ID>DATA_OUT_1</ID>129 </output>
<output>
<ID>DATA_OUT_2</ID>125 </output>
<output>
<ID>DATA_OUT_3</ID>124 </output>
<output>
<ID>DATA_OUT_4</ID>123 </output>
<output>
<ID>DATA_OUT_5</ID>121 </output>
<output>
<ID>DATA_OUT_6</ID>120 </output>
<output>
<ID>DATA_OUT_7</ID>119 </output>
<input>
<ID>ENABLE_0</ID>197 </input>
<input>
<ID>write_clock</ID>193 </input>
<input>
<ID>write_enable</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 121</lparam>
<lparam>Address:1 113</lparam>
<lparam>Address:2 123</lparam>
<lparam>Address:3 117</lparam>
<lparam>Address:4 108</lparam>
<lparam>Address:5 106</lparam>
<lparam>Address:13 4</lparam></gate>
<gate>
<ID>112</ID>
<type>EE_VDD</type>
<position>-210,5.5</position>
<output>
<ID>OUT_0</ID>197 </output>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>114</ID>
<type>DE_TO</type>
<position>-185,-17.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-REG-IN</lparam></gate>
<gate>
<ID>505</ID>
<type>DA_FROM</type>
<position>-238,33</position>
<input>
<ID>IN_0</ID>433 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-IN-1</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>-194,6</position>
<input>
<ID>IN_0</ID>378 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID READY-TO-SAVE-INSTRUCTION</lparam></gate>
<gate>
<ID>508</ID>
<type>DA_FROM</type>
<position>-238,38</position>
<input>
<ID>IN_0</ID>432 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-IN-2</lparam></gate>
<gate>
<ID>510</ID>
<type>DA_FROM</type>
<position>-238,43</position>
<input>
<ID>IN_0</ID>431 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID MBR-IN-3</lparam></gate>
<gate>
<ID>511</ID>
<type>AA_MUX_2x1</type>
<position>-225,57</position>
<input>
<ID>IN_0</ID>549 </input>
<input>
<ID>IN_1</ID>427 </input>
<output>
<ID>OUT</ID>419 </output>
<input>
<ID>SEL_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>512</ID>
<type>DA_FROM</type>
<position>-235.5,85</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-3</lparam></gate>
<gate>
<ID>513</ID>
<type>DA_FROM</type>
<position>-235.5,77.5</position>
<input>
<ID>IN_0</ID>420 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-0</lparam></gate>
<gate>
<ID>900</ID>
<type>AE_OR2</type>
<position>-209,9.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>639 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_LABEL</type>
<position>-210.5,17.5</position>
<gparam>LABEL_TEXT 16 x 8-bit Instruction RAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>516</ID>
<type>DA_FROM</type>
<position>-235.5,80</position>
<input>
<ID>IN_0</ID>558 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-1</lparam></gate>
<gate>
<ID>130</ID>
<type>DE_TO</type>
<position>-185,-21.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-3-IN</lparam></gate>
<gate>
<ID>517</ID>
<type>AA_MUX_2x1</type>
<position>-225,52</position>
<input>
<ID>IN_0</ID>550 </input>
<input>
<ID>IN_1</ID>428 </input>
<output>
<ID>OUT</ID>421 </output>
<input>
<ID>SEL_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>518</ID>
<type>AA_MUX_2x1</type>
<position>-225,47</position>
<input>
<ID>IN_0</ID>551 </input>
<input>
<ID>IN_1</ID>430 </input>
<output>
<ID>OUT</ID>422 </output>
<input>
<ID>SEL_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>DE_TO</type>
<position>-185,-25.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-2-IN</lparam></gate>
<gate>
<ID>519</ID>
<type>GA_LED</type>
<position>-186.5,76.5</position>
<input>
<ID>N_in0</ID>434 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>520</ID>
<type>AA_MUX_2x1</type>
<position>-225,42</position>
<input>
<ID>IN_0</ID>552 </input>
<input>
<ID>IN_1</ID>431 </input>
<output>
<ID>OUT</ID>423 </output>
<input>
<ID>SEL_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AA_LABEL</type>
<position>-245,-10.5</position>
<gparam>LABEL_TEXT Input Instruction</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>522</ID>
<type>DA_FROM</type>
<position>-215.5,53</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID LOAD-MBR</lparam></gate>
<gate>
<ID>336</ID>
<type>AA_AND2</type>
<position>-199,7</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>530 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>-185,-29.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-1-IN</lparam></gate>
<gate>
<ID>338</ID>
<type>AA_MUX_2x1</type>
<position>-227.5,-19.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>619 </input>
<output>
<ID>OUT</ID>113 </output>
<input>
<ID>SEL_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>DE_TO</type>
<position>-185,-33.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-0-IN</lparam></gate>
<gate>
<ID>147</ID>
<type>DE_TO</type>
<position>-185,-37.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-2-IN</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>-185,-41.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-1-IN</lparam></gate>
<gate>
<ID>351</ID>
<type>DA_FROM</type>
<position>-238,8.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-RAM-3</lparam></gate>
<gate>
<ID>545</ID>
<type>AA_MUX_2x1</type>
<position>-225,37</position>
<input>
<ID>IN_0</ID>557 </input>
<input>
<ID>IN_1</ID>432 </input>
<output>
<ID>OUT</ID>424 </output>
<input>
<ID>SEL_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>DA_FROM</type>
<position>-238,1</position>
<input>
<ID>IN_0</ID>669 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-RAM-0</lparam></gate>
<gate>
<ID>546</ID>
<type>AA_MUX_2x1</type>
<position>-225,32</position>
<input>
<ID>IN_0</ID>560 </input>
<input>
<ID>IN_1</ID>433 </input>
<output>
<ID>OUT</ID>425 </output>
<input>
<ID>SEL_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>DA_FROM</type>
<position>-238,3.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-RAM-1</lparam></gate>
<gate>
<ID>547</ID>
<type>AA_TOGGLE</type>
<position>-208.5,37</position>
<output>
<ID>OUT_0</ID>579 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_MUX_2x1</type>
<position>-227.5,-24.5</position>
<input>
<ID>IN_0</ID>121 </input>
<input>
<ID>IN_1</ID>620 </input>
<output>
<ID>OUT</ID>114 </output>
<input>
<ID>SEL_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_MUX_2x1</type>
<position>-227.5,-29.5</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>621 </input>
<output>
<ID>OUT</ID>115 </output>
<input>
<ID>SEL_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>DA_FROM</type>
<position>-233.5,-1.5</position>
<input>
<ID>IN_0</ID>541 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID USE-USER-INSTRUCTION</lparam></gate>
<gate>
<ID>365</ID>
<type>AA_MUX_2x1</type>
<position>-227.5,-34.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>622 </input>
<output>
<ID>OUT</ID>116 </output>
<input>
<ID>SEL_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>385</ID>
<type>AA_MUX_2x1</type>
<position>-227.5,-39.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>623 </input>
<output>
<ID>OUT</ID>117 </output>
<input>
<ID>SEL_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>26</ID>
<points>-214.5,6,-214.5,9.5</points>
<connection>
<GID>111</GID>
<name>write_clock</name></connection>
<intersection>9.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>-214.5,9.5,-212,9.5</points>
<connection>
<GID>900</GID>
<name>OUT</name></connection>
<intersection>-214.5 26</intersection></hsegment></shape></wire>
<wire>
<ID>579</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-208.5,39,-208.5,40</points>
<connection>
<GID>547</GID>
<name>OUT_0</name></connection>
<intersection>40 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-210,40,-208.5,40</points>
<connection>
<GID>460</GID>
<name>clear</name></connection>
<intersection>-208.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-226.5,5,-226.5,13.5</points>
<intersection>5 6</intersection>
<intersection>7 4</intersection>
<intersection>8 1</intersection>
<intersection>13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-226.5,8,-224.5,8</points>
<connection>
<GID>111</GID>
<name>ADDRESS_7</name></connection>
<intersection>-226.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-235,13.5,-226.5,13.5</points>
<intersection>-235 9</intersection>
<intersection>-226.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-226.5,7,-224.5,7</points>
<connection>
<GID>111</GID>
<name>ADDRESS_6</name></connection>
<intersection>-226.5 0</intersection>
<intersection>-224.5 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-226.5,5,-224.5,5</points>
<connection>
<GID>111</GID>
<name>ADDRESS_4</name></connection>
<intersection>-226.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-224.5,6,-224.5,7</points>
<connection>
<GID>111</GID>
<name>ADDRESS_5</name></connection>
<intersection>7 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-235,12.5,-235,13.5</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>13.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-215.5,51,-212,51</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<connection>
<GID>460</GID>
<name>load</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-214.5,4,-210,4</points>
<connection>
<GID>111</GID>
<name>ENABLE_0</name></connection>
<intersection>-210 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-210,4,-210,4.5</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>4 1</intersection></vsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-189.5,-49.5,-189.5,-12.5</points>
<connection>
<GID>76</GID>
<name>T_in2</name></connection>
<intersection>-49.5 10</intersection>
<intersection>-45.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-189.5,-45.5,-187,-45.5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>-189.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-225.5,-49.5,-189.5,-49.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>-189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>417</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,63,-227,63</points>
<connection>
<GID>473</GID>
<name>IN_1</name></connection>
<connection>
<GID>458</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-217,49,-217,62</points>
<intersection>49 6</intersection>
<intersection>62 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-223,62,-217,62</points>
<connection>
<GID>473</GID>
<name>OUT</name></connection>
<intersection>-217 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-217,49,-215,49</points>
<connection>
<GID>460</GID>
<name>IN_7</name></connection>
<intersection>-217 0</intersection></hsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-218,48,-218,57</points>
<intersection>48 1</intersection>
<intersection>57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-218,48,-215,48</points>
<connection>
<GID>460</GID>
<name>IN_6</name></connection>
<intersection>-218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-223,57,-218,57</points>
<connection>
<GID>511</GID>
<name>OUT</name></connection>
<intersection>-218 0</intersection></hsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-233.5,77.5,-222,77.5</points>
<connection>
<GID>679</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>513</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-220,47,-220,52</points>
<intersection>47 1</intersection>
<intersection>52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-220,47,-215,47</points>
<connection>
<GID>460</GID>
<name>IN_5</name></connection>
<intersection>-220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-223,52,-220,52</points>
<connection>
<GID>517</GID>
<name>OUT</name></connection>
<intersection>-220 0</intersection></hsegment></shape></wire>
<wire>
<ID>422</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-223,46,-215,46</points>
<connection>
<GID>460</GID>
<name>IN_4</name></connection>
<intersection>-223 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-223,46,-223,47</points>
<connection>
<GID>518</GID>
<name>OUT</name></connection>
<intersection>46 1</intersection></vsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-219,42,-219,45</points>
<intersection>42 2</intersection>
<intersection>45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-219,45,-215,45</points>
<connection>
<GID>460</GID>
<name>IN_3</name></connection>
<intersection>-219 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-223,42,-219,42</points>
<connection>
<GID>520</GID>
<name>OUT</name></connection>
<intersection>-219 0</intersection></hsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-218,37,-218,44</points>
<intersection>37 2</intersection>
<intersection>44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-218,44,-215,44</points>
<connection>
<GID>460</GID>
<name>IN_2</name></connection>
<intersection>-218 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-223,37,-218,37</points>
<connection>
<GID>545</GID>
<name>OUT</name></connection>
<intersection>-218 0</intersection></hsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-217,32,-217,43</points>
<intersection>32 2</intersection>
<intersection>43 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-217,43,-215,43</points>
<connection>
<GID>460</GID>
<name>IN_1</name></connection>
<intersection>-217 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-223,32,-217,32</points>
<connection>
<GID>546</GID>
<name>OUT</name></connection>
<intersection>-217 0</intersection></hsegment></shape></wire>
<wire>
<ID>618</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239.5,-13.5,-229.5,-13.5</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<connection>
<GID>826</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>619</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-18.5,-229.5,-18.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<connection>
<GID>827</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-216,27,-216,42</points>
<intersection>27 2</intersection>
<intersection>42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-216,42,-215,42</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>-216 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-223,27,-216,27</points>
<connection>
<GID>629</GID>
<name>OUT</name></connection>
<intersection>-216 0</intersection></hsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,58,-227,58</points>
<connection>
<GID>511</GID>
<name>IN_1</name></connection>
<connection>
<GID>457</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>620</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-23.5,-229.5,-23.5</points>
<connection>
<GID>354</GID>
<name>IN_1</name></connection>
<connection>
<GID>829</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,53,-227,53</points>
<connection>
<GID>517</GID>
<name>IN_1</name></connection>
<connection>
<GID>454</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>621</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-28.5,-229.5,-28.5</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<connection>
<GID>830</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>622</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-33.5,-229.5,-33.5</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<connection>
<GID>832</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,48,-227,48</points>
<connection>
<GID>518</GID>
<name>IN_1</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>623</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-38.5,-229.5,-38.5</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<connection>
<GID>385</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,43,-227,43</points>
<connection>
<GID>520</GID>
<name>IN_1</name></connection>
<connection>
<GID>510</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>624</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-48.5,-229.5,-48.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<connection>
<GID>835</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,38,-227,38</points>
<connection>
<GID>545</GID>
<name>IN_1</name></connection>
<connection>
<GID>508</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>625</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-239,-43.5,-229.5,-43.5</points>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<connection>
<GID>834</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,33,-227,33</points>
<connection>
<GID>546</GID>
<name>IN_1</name></connection>
<connection>
<GID>505</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-222,74,-188,74</points>
<intersection>-222 90</intersection>
<intersection>-209 19</intersection>
<intersection>-206 112</intersection>
<intersection>-203 107</intersection>
<intersection>-200 108</intersection>
<intersection>-197 109</intersection>
<intersection>-194 110</intersection>
<intersection>-191 111</intersection>
<intersection>-188 113</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-209,67,-209,81.5</points>
<connection>
<GID>464</GID>
<name>T_ctrl</name></connection>
<intersection>74 1</intersection>
<intersection>81.5 48</intersection></vsegment>
<hsegment>
<ID>48</ID>
<points>-212,81.5,-209,81.5</points>
<connection>
<GID>679</GID>
<name>write_enable</name></connection>
<intersection>-209 19</intersection></hsegment>
<vsegment>
<ID>90</ID>
<points>-222,29.5,-222,74</points>
<intersection>29.5 92</intersection>
<intersection>34.5 99</intersection>
<intersection>39.5 98</intersection>
<intersection>44.5 97</intersection>
<intersection>49.5 96</intersection>
<intersection>54.5 95</intersection>
<intersection>59.5 94</intersection>
<intersection>64.5 93</intersection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>92</ID>
<points>-225,29.5,-222,29.5</points>
<connection>
<GID>629</GID>
<name>SEL_0</name></connection>
<intersection>-222 90</intersection></hsegment>
<hsegment>
<ID>93</ID>
<points>-225,64.5,-222,64.5</points>
<connection>
<GID>473</GID>
<name>SEL_0</name></connection>
<intersection>-222 90</intersection></hsegment>
<hsegment>
<ID>94</ID>
<points>-225,59.5,-222,59.5</points>
<connection>
<GID>511</GID>
<name>SEL_0</name></connection>
<intersection>-222 90</intersection></hsegment>
<hsegment>
<ID>95</ID>
<points>-225,54.5,-222,54.5</points>
<connection>
<GID>517</GID>
<name>SEL_0</name></connection>
<intersection>-222 90</intersection></hsegment>
<hsegment>
<ID>96</ID>
<points>-225,49.5,-222,49.5</points>
<connection>
<GID>518</GID>
<name>SEL_0</name></connection>
<intersection>-222 90</intersection></hsegment>
<hsegment>
<ID>97</ID>
<points>-225,44.5,-222,44.5</points>
<connection>
<GID>520</GID>
<name>SEL_0</name></connection>
<intersection>-222 90</intersection></hsegment>
<hsegment>
<ID>98</ID>
<points>-225,39.5,-222,39.5</points>
<connection>
<GID>545</GID>
<name>SEL_0</name></connection>
<intersection>-222 90</intersection></hsegment>
<hsegment>
<ID>99</ID>
<points>-225,34.5,-222,34.5</points>
<connection>
<GID>546</GID>
<name>SEL_0</name></connection>
<intersection>-222 90</intersection></hsegment>
<vsegment>
<ID>107</ID>
<points>-203,67,-203,74</points>
<connection>
<GID>632</GID>
<name>T_ctrl</name></connection>
<intersection>74 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-200,67,-200,74</points>
<connection>
<GID>633</GID>
<name>T_ctrl</name></connection>
<intersection>74 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-197,67,-197,74</points>
<connection>
<GID>634</GID>
<name>T_ctrl</name></connection>
<intersection>74 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-194,67,-194,74</points>
<connection>
<GID>635</GID>
<name>T_ctrl</name></connection>
<intersection>74 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-191,67,-191,79.5</points>
<connection>
<GID>636</GID>
<name>T_ctrl</name></connection>
<intersection>74 1</intersection>
<intersection>76.5 130</intersection>
<intersection>79.5 127</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>-206,67,-206,74</points>
<connection>
<GID>630</GID>
<name>T_ctrl</name></connection>
<intersection>74 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>-188,67,-188,74</points>
<connection>
<GID>638</GID>
<name>T_ctrl</name></connection>
<intersection>74 1</intersection></vsegment>
<hsegment>
<ID>127</ID>
<points>-191,79.5,-190,79.5</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>-191 111</intersection></hsegment>
<hsegment>
<ID>130</ID>
<points>-191,76.5,-187.5,76.5</points>
<connection>
<GID>519</GID>
<name>N_in0</name></connection>
<intersection>-191 111</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,28,-227,28</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<connection>
<GID>629</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-207,49,-207,63</points>
<connection>
<GID>460</GID>
<name>OUT_7</name></connection>
<intersection>59 1</intersection>
<intersection>63 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-207,59,-184.5,59</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<intersection>-207 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-208,63,-207,63</points>
<intersection>-208 3</intersection>
<intersection>-207 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-208,63,-208,64</points>
<connection>
<GID>464</GID>
<name>T_in2</name></connection>
<intersection>63 2</intersection></vsegment></shape></wire>
<wire>
<ID>639</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-206,10.5,-204,10.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>-206 1</intersection></hsegment>
<vsegment>
<ID>1</ID>
<points>-206,10.5,-206,10.5</points>
<connection>
<GID>900</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection></vsegment></shape></wire>
<wire>
<ID>669</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-236,1,-224.5,1</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>ADDRESS_0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-213.5,-2.5,-190.5,-2.5</points>
<intersection>-213.5 151</intersection>
<intersection>-211.5 148</intersection>
<intersection>-208.5 112</intersection>
<intersection>-205.5 107</intersection>
<intersection>-204 19</intersection>
<intersection>-202.5 108</intersection>
<intersection>-199.5 109</intersection>
<intersection>-196.5 110</intersection>
<intersection>-193.5 111</intersection>
<intersection>-190.5 113</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-204,-2.5,-204,8.5</points>
<intersection>-2.5 1</intersection>
<intersection>7 154</intersection>
<intersection>8.5 152</intersection></vsegment>
<vsegment>
<ID>107</ID>
<points>-205.5,-9.5,-205.5,-2.5</points>
<connection>
<GID>67</GID>
<name>T_ctrl</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>108</ID>
<points>-202.5,-9.5,-202.5,-2.5</points>
<connection>
<GID>69</GID>
<name>T_ctrl</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>109</ID>
<points>-199.5,-9.5,-199.5,-2.5</points>
<connection>
<GID>70</GID>
<name>T_ctrl</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>110</ID>
<points>-196.5,-9.5,-196.5,-2.5</points>
<connection>
<GID>71</GID>
<name>T_ctrl</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>111</ID>
<points>-193.5,-9.5,-193.5,-2.5</points>
<connection>
<GID>75</GID>
<name>T_ctrl</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>112</ID>
<points>-208.5,-9.5,-208.5,-2.5</points>
<connection>
<GID>65</GID>
<name>T_ctrl</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>-190.5,-9.5,-190.5,-2.5</points>
<connection>
<GID>76</GID>
<name>T_ctrl</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>148</ID>
<points>-211.5,-9.5,-211.5,-2.5</points>
<connection>
<GID>98</GID>
<name>T_ctrl</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>151</ID>
<points>-213.5,-2.5,-213.5,5</points>
<intersection>-2.5 1</intersection>
<intersection>5 153</intersection></vsegment>
<hsegment>
<ID>152</ID>
<points>-206,8.5,-204,8.5</points>
<connection>
<GID>900</GID>
<name>IN_0</name></connection>
<intersection>-204 19</intersection></hsegment>
<hsegment>
<ID>153</ID>
<points>-214.5,5,-213.5,5</points>
<connection>
<GID>111</GID>
<name>write_enable</name></connection>
<intersection>-213.5 151</intersection></hsegment>
<hsegment>
<ID>154</ID>
<points>-204,7,-202,7</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<intersection>-204 19</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-210.5,-17.5,-210.5,-12.5</points>
<connection>
<GID>98</GID>
<name>T_in2</name></connection>
<intersection>-17.5 6</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-225.5,-14.5,-210.5,-14.5</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>-210.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-210.5,-17.5,-187,-17.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-210.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-207.5,-21.5,-207.5,-12.5</points>
<connection>
<GID>65</GID>
<name>T_in2</name></connection>
<intersection>-21.5 7</intersection>
<intersection>-19.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-207.5,-21.5,-187,-21.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-207.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-225.5,-19.5,-207.5,-19.5</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>-207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-204.5,-25.5,-204.5,-12.5</points>
<connection>
<GID>67</GID>
<name>T_in2</name></connection>
<intersection>-25.5 7</intersection>
<intersection>-24.5 9</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-204.5,-25.5,-187,-25.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-204.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-225.5,-24.5,-204.5,-24.5</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<intersection>-204.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-201.5,-29.5,-201.5,-12.5</points>
<connection>
<GID>69</GID>
<name>T_in2</name></connection>
<intersection>-29.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-225.5,-29.5,-187,-29.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<intersection>-201.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-198.5,-34.5,-198.5,-12.5</points>
<connection>
<GID>70</GID>
<name>T_in2</name></connection>
<intersection>-34.5 8</intersection>
<intersection>-33.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-198.5,-33.5,-187,-33.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-198.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-225.5,-34.5,-198.5,-34.5</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<intersection>-198.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-195.5,-39.5,-195.5,-12.5</points>
<connection>
<GID>71</GID>
<name>T_in2</name></connection>
<intersection>-39.5 8</intersection>
<intersection>-37.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-195.5,-37.5,-187,-37.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>-195.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-225.5,-39.5,-195.5,-39.5</points>
<connection>
<GID>385</GID>
<name>OUT</name></connection>
<intersection>-195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-192.5,-44.5,-192.5,-12.5</points>
<connection>
<GID>75</GID>
<name>T_in2</name></connection>
<intersection>-44.5 8</intersection>
<intersection>-41.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-192.5,-41.5,-187,-41.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-192.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-225.5,-44.5,-192.5,-44.5</points>
<connection>
<GID>389</GID>
<name>OUT</name></connection>
<intersection>-192.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230.5,-15.5,-230.5,-11</points>
<intersection>-15.5 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-230.5,-15.5,-229.5,-15.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>-230.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-230.5,-11,-214,-11</points>
<intersection>-230.5 0</intersection>
<intersection>-223 3</intersection>
<intersection>-214 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-223,-11,-223,-2.5</points>
<connection>
<GID>111</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>111</GID>
<name>DATA_IN_7</name></connection>
<intersection>-11 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-214,-12.5,-214,-11</points>
<intersection>-12.5 5</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-214,-12.5,-212.5,-12.5</points>
<connection>
<GID>98</GID>
<name>T_in</name></connection>
<intersection>-214 4</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-231.5,-20.5,-231.5,-10</points>
<intersection>-20.5 1</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-231.5,-20.5,-229.5,-20.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>-231.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-231.5,-10,-210,-10</points>
<intersection>-231.5 0</intersection>
<intersection>-222 3</intersection>
<intersection>-210 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-222,-10,-222,-2.5</points>
<connection>
<GID>111</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>111</GID>
<name>DATA_IN_6</name></connection>
<intersection>-10 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-210,-12.5,-210,-10</points>
<intersection>-12.5 5</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-210,-12.5,-209.5,-12.5</points>
<connection>
<GID>65</GID>
<name>T_in</name></connection>
<intersection>-210 4</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-232.5,-25.5,-232.5,-8</points>
<intersection>-25.5 1</intersection>
<intersection>-8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-232.5,-25.5,-229.5,-25.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>-232.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-232.5,-8,-206.5,-8</points>
<intersection>-232.5 0</intersection>
<intersection>-221 3</intersection>
<intersection>-206.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-221,-8,-221,-2.5</points>
<connection>
<GID>111</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>111</GID>
<name>DATA_IN_5</name></connection>
<intersection>-8 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-206.5,-12.5,-206.5,-8</points>
<connection>
<GID>67</GID>
<name>T_in</name></connection>
<intersection>-8 2</intersection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-233.5,-30.5,-233.5,-9</points>
<intersection>-30.5 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233.5,-30.5,-229.5,-30.5</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>-233.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233.5,-9,-203.5,-9</points>
<intersection>-233.5 0</intersection>
<intersection>-220 3</intersection>
<intersection>-203.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-220,-9,-220,-2.5</points>
<connection>
<GID>111</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>111</GID>
<name>DATA_IN_4</name></connection>
<intersection>-9 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-203.5,-12.5,-203.5,-9</points>
<connection>
<GID>69</GID>
<name>T_in</name></connection>
<intersection>-9 2</intersection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-234.5,-35.5,-234.5,-7</points>
<intersection>-35.5 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-234.5,-35.5,-229.5,-35.5</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>-234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-234.5,-7,-200.5,-7</points>
<intersection>-234.5 0</intersection>
<intersection>-219 3</intersection>
<intersection>-200.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-219,-7,-219,-2.5</points>
<connection>
<GID>111</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>111</GID>
<name>DATA_IN_3</name></connection>
<intersection>-7 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-200.5,-12.5,-200.5,-7</points>
<connection>
<GID>70</GID>
<name>T_in</name></connection>
<intersection>-7 2</intersection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-235.5,-40.5,-235.5,-6</points>
<intersection>-40.5 1</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-235.5,-40.5,-229.5,-40.5</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>-235.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-235.5,-6,-197.5,-6</points>
<intersection>-235.5 0</intersection>
<intersection>-218 3</intersection>
<intersection>-197.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-218,-6,-218,-2.5</points>
<connection>
<GID>111</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>111</GID>
<name>DATA_IN_2</name></connection>
<intersection>-6 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-197.5,-12.5,-197.5,-6</points>
<connection>
<GID>71</GID>
<name>T_in</name></connection>
<intersection>-6 2</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-234.5,2,-234.5,3.5</points>
<intersection>2 1</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-234.5,2,-224.5,2</points>
<connection>
<GID>111</GID>
<name>ADDRESS_1</name></connection>
<intersection>-234.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-236,3.5,-234.5,3.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-236.5,-45.5,-236.5,-5</points>
<intersection>-45.5 1</intersection>
<intersection>-5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-236.5,-45.5,-229.5,-45.5</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-236.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-236.5,-5,-194.5,-5</points>
<intersection>-236.5 0</intersection>
<intersection>-217 3</intersection>
<intersection>-194.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-217,-5,-217,-2.5</points>
<connection>
<GID>111</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>111</GID>
<name>DATA_IN_1</name></connection>
<intersection>-5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-194.5,-12.5,-194.5,-5</points>
<connection>
<GID>75</GID>
<name>T_in</name></connection>
<intersection>-5 2</intersection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-237.5,-50.5,-237.5,-3.5</points>
<intersection>-50.5 1</intersection>
<intersection>-3.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-237.5,-50.5,-229.5,-50.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-237.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-237.5,-3.5,-191.5,-3.5</points>
<intersection>-237.5 0</intersection>
<intersection>-216 4</intersection>
<intersection>-191.5 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-216,-3.5,-216,-2.5</points>
<connection>
<GID>111</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>111</GID>
<name>DATA_IN_0</name></connection>
<intersection>-3.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-191.5,-12.5,-191.5,-3.5</points>
<connection>
<GID>76</GID>
<name>T_in</name></connection>
<intersection>-3.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-233.5,3,-233.5,6</points>
<intersection>3 1</intersection>
<intersection>6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233.5,3,-224.5,3</points>
<connection>
<GID>111</GID>
<name>ADDRESS_2</name></connection>
<intersection>-233.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-236,6,-233.5,6</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-233.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>530</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-196,8,-196,8</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>336</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230.5,4,-230.5,8.5</points>
<intersection>4 1</intersection>
<intersection>8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-230.5,4,-224.5,4</points>
<connection>
<GID>111</GID>
<name>ADDRESS_3</name></connection>
<intersection>-230.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-236,8.5,-230.5,8.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-230.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>541</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-224.5,-47,-224.5,-1.5</points>
<intersection>-47 9</intersection>
<intersection>-42 10</intersection>
<intersection>-37 11</intersection>
<intersection>-32 12</intersection>
<intersection>-27 13</intersection>
<intersection>-22 14</intersection>
<intersection>-17 15</intersection>
<intersection>-12 58</intersection>
<intersection>-1.5 60</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-227.5,-47,-224.5,-47</points>
<connection>
<GID>62</GID>
<name>SEL_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-227.5,-42,-224.5,-42</points>
<connection>
<GID>389</GID>
<name>SEL_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-227.5,-37,-224.5,-37</points>
<connection>
<GID>385</GID>
<name>SEL_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-227.5,-32,-224.5,-32</points>
<connection>
<GID>365</GID>
<name>SEL_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-227.5,-27,-224.5,-27</points>
<connection>
<GID>363</GID>
<name>SEL_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-227.5,-22,-224.5,-22</points>
<connection>
<GID>354</GID>
<name>SEL_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-227.5,-17,-224.5,-17</points>
<connection>
<GID>338</GID>
<name>SEL_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>58</ID>
<points>-227.5,-12,-224.5,-12</points>
<connection>
<GID>99</GID>
<name>SEL_0</name></connection>
<intersection>-224.5 0</intersection></hsegment>
<hsegment>
<ID>60</ID>
<points>-231.5,-1.5,-224.5,-1.5</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-224.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>542</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-206,48,-206,63</points>
<intersection>48 2</intersection>
<intersection>55 1</intersection>
<intersection>63 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-206,55,-184.5,55</points>
<connection>
<GID>682</GID>
<name>IN_0</name></connection>
<intersection>-206 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-207,48,-206,48</points>
<connection>
<GID>460</GID>
<name>OUT_6</name></connection>
<intersection>-206 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-206,63,-205,63</points>
<intersection>-206 0</intersection>
<intersection>-205 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-205,63,-205,64</points>
<connection>
<GID>630</GID>
<name>T_in2</name></connection>
<intersection>63 4</intersection></vsegment></shape></wire>
<wire>
<ID>543</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-205,47,-205,62</points>
<intersection>47 1</intersection>
<intersection>51 2</intersection>
<intersection>62 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-207,47,-205,47</points>
<connection>
<GID>460</GID>
<name>OUT_5</name></connection>
<intersection>-205 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-205,51,-184.5,51</points>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>-205 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-205,62,-202,62</points>
<intersection>-205 0</intersection>
<intersection>-202 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-202,62,-202,64</points>
<connection>
<GID>632</GID>
<name>T_in2</name></connection>
<intersection>62 4</intersection></vsegment></shape></wire>
<wire>
<ID>544</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-207,46,-184.5,46</points>
<connection>
<GID>460</GID>
<name>OUT_4</name></connection>
<intersection>-204 2</intersection>
<intersection>-184.5 5</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-204,46,-204,61.5</points>
<intersection>46 1</intersection>
<intersection>61.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-204,61.5,-199,61.5</points>
<intersection>-204 2</intersection>
<intersection>-199 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-199,61.5,-199,64</points>
<connection>
<GID>633</GID>
<name>T_in2</name></connection>
<intersection>61.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-184.5,46,-184.5,47</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<intersection>46 1</intersection></vsegment></shape></wire>
<wire>
<ID>545</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-201,43,-201,61</points>
<intersection>43 1</intersection>
<intersection>45 2</intersection>
<intersection>61 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-201,43,-184.5,43</points>
<connection>
<GID>685</GID>
<name>IN_0</name></connection>
<intersection>-201 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-207,45,-201,45</points>
<connection>
<GID>460</GID>
<name>OUT_3</name></connection>
<intersection>-201 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-201,61,-196,61</points>
<intersection>-201 0</intersection>
<intersection>-196 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-196,61,-196,64</points>
<connection>
<GID>634</GID>
<name>T_in2</name></connection>
<intersection>61 3</intersection></vsegment></shape></wire>
<wire>
<ID>546</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-200,39,-200,60.5</points>
<intersection>39 1</intersection>
<intersection>44 2</intersection>
<intersection>60.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-200,39,-184.5,39</points>
<connection>
<GID>686</GID>
<name>IN_0</name></connection>
<intersection>-200 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-207,44,-200,44</points>
<connection>
<GID>460</GID>
<name>OUT_2</name></connection>
<intersection>-200 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-200,60.5,-193,60.5</points>
<intersection>-200 0</intersection>
<intersection>-193 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-193,60.5,-193,64</points>
<connection>
<GID>635</GID>
<name>T_in2</name></connection>
<intersection>60.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>547</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-199,35,-199,60</points>
<intersection>35 2</intersection>
<intersection>43 1</intersection>
<intersection>60 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-207,43,-199,43</points>
<connection>
<GID>460</GID>
<name>OUT_1</name></connection>
<intersection>-199 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-199,35,-184.5,35</points>
<connection>
<GID>687</GID>
<name>IN_0</name></connection>
<intersection>-199 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-199,60,-190,60</points>
<intersection>-199 0</intersection>
<intersection>-190 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-190,60,-190,64</points>
<connection>
<GID>636</GID>
<name>T_in2</name></connection>
<intersection>60 3</intersection></vsegment></shape></wire>
<wire>
<ID>548</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-228,61,-228,65.5</points>
<intersection>61 1</intersection>
<intersection>65.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-228,61,-227,61</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>-228 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-228,65.5,-211.5,65.5</points>
<intersection>-228 0</intersection>
<intersection>-220.5 3</intersection>
<intersection>-211.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-220.5,65.5,-220.5,74</points>
<connection>
<GID>679</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>679</GID>
<name>DATA_IN_7</name></connection>
<intersection>65.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-211.5,64,-211.5,65.5</points>
<intersection>64 5</intersection>
<intersection>65.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-211.5,64,-210,64</points>
<connection>
<GID>464</GID>
<name>T_in</name></connection>
<intersection>-211.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>549</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-229,56,-229,66.5</points>
<intersection>56 1</intersection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-229,56,-227,56</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<intersection>-229 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-229,66.5,-207.5,66.5</points>
<intersection>-229 0</intersection>
<intersection>-219.5 3</intersection>
<intersection>-207.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-219.5,66.5,-219.5,74</points>
<connection>
<GID>679</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>679</GID>
<name>DATA_IN_6</name></connection>
<intersection>66.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-207.5,64,-207.5,66.5</points>
<intersection>64 5</intersection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-207.5,64,-207,64</points>
<connection>
<GID>630</GID>
<name>T_in</name></connection>
<intersection>-207.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>550</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-230,51,-230,67.5</points>
<intersection>51 1</intersection>
<intersection>67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-230,51,-227,51</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<intersection>-230 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-230,67.5,-204,67.5</points>
<intersection>-230 0</intersection>
<intersection>-218.5 3</intersection>
<intersection>-204 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-218.5,67.5,-218.5,74</points>
<connection>
<GID>679</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>679</GID>
<name>DATA_IN_5</name></connection>
<intersection>67.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-204,64,-204,67.5</points>
<connection>
<GID>632</GID>
<name>T_in</name></connection>
<intersection>67.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>551</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-231,46,-231,68.5</points>
<intersection>46 1</intersection>
<intersection>68.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-231,46,-227,46</points>
<connection>
<GID>518</GID>
<name>IN_0</name></connection>
<intersection>-231 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-231,68.5,-201,68.5</points>
<intersection>-231 0</intersection>
<intersection>-217.5 3</intersection>
<intersection>-201 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-217.5,68.5,-217.5,74</points>
<connection>
<GID>679</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>679</GID>
<name>DATA_IN_4</name></connection>
<intersection>68.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-201,64,-201,68.5</points>
<connection>
<GID>633</GID>
<name>T_in</name></connection>
<intersection>68.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>552</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-232,41,-232,69.5</points>
<intersection>41 1</intersection>
<intersection>69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-232,41,-227,41</points>
<connection>
<GID>520</GID>
<name>IN_0</name></connection>
<intersection>-232 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-232,69.5,-198,69.5</points>
<intersection>-232 0</intersection>
<intersection>-216.5 3</intersection>
<intersection>-198 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-216.5,69.5,-216.5,74</points>
<connection>
<GID>679</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>679</GID>
<name>DATA_IN_3</name></connection>
<intersection>69.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-198,64,-198,69.5</points>
<connection>
<GID>634</GID>
<name>T_in</name></connection>
<intersection>69.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>557</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-233,36,-233,70.5</points>
<intersection>36 1</intersection>
<intersection>70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-233,36,-227,36</points>
<connection>
<GID>545</GID>
<name>IN_0</name></connection>
<intersection>-233 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233,70.5,-195,70.5</points>
<intersection>-233 0</intersection>
<intersection>-215.5 3</intersection>
<intersection>-195 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-215.5,70.5,-215.5,74</points>
<connection>
<GID>679</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>679</GID>
<name>DATA_IN_2</name></connection>
<intersection>70.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-195,64,-195,70.5</points>
<connection>
<GID>635</GID>
<name>T_in</name></connection>
<intersection>70.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>558</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-232,78.5,-232,80</points>
<intersection>78.5 1</intersection>
<intersection>80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-232,78.5,-222,78.5</points>
<connection>
<GID>679</GID>
<name>ADDRESS_1</name></connection>
<intersection>-232 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233.5,80,-232,80</points>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>-232 0</intersection></hsegment></shape></wire>
<wire>
<ID>560</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-234,31,-234,71.5</points>
<intersection>31 1</intersection>
<intersection>71.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-234,31,-227,31</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<intersection>-234 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-234,71.5,-192,71.5</points>
<intersection>-234 0</intersection>
<intersection>-214.5 3</intersection>
<intersection>-192 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-214.5,71.5,-214.5,74</points>
<connection>
<GID>679</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>679</GID>
<name>DATA_IN_1</name></connection>
<intersection>71.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-192,64,-192,71.5</points>
<connection>
<GID>636</GID>
<name>T_in</name></connection>
<intersection>71.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>568</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-235,26,-235,73</points>
<intersection>26 1</intersection>
<intersection>73 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-235,26,-227,26</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<intersection>-235 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-235,73,-189,73</points>
<intersection>-235 0</intersection>
<intersection>-213.5 4</intersection>
<intersection>-189 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-213.5,73,-213.5,74</points>
<connection>
<GID>679</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>679</GID>
<name>DATA_IN_0</name></connection>
<intersection>73 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-189,64,-189,73</points>
<connection>
<GID>638</GID>
<name>T_in</name></connection>
<intersection>73 3</intersection></vsegment></shape></wire>
<wire>
<ID>569</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-231,79.5,-231,82.5</points>
<intersection>79.5 1</intersection>
<intersection>82.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-231,79.5,-222,79.5</points>
<connection>
<GID>679</GID>
<name>ADDRESS_2</name></connection>
<intersection>-231 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233.5,82.5,-231,82.5</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<intersection>-231 0</intersection></hsegment></shape></wire>
<wire>
<ID>570</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-228,80.5,-228,85</points>
<intersection>80.5 1</intersection>
<intersection>85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-228,80.5,-222,80.5</points>
<connection>
<GID>679</GID>
<name>ADDRESS_3</name></connection>
<intersection>-228 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-233.5,85,-228,85</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<intersection>-228 0</intersection></hsegment></shape></wire>
<wire>
<ID>378</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-196,6,-196,6</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-196,6,-196,6</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-196 0</intersection></hsegment></shape></wire>
<wire>
<ID>572</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-212,82.5,-167.5,82.5</points>
<connection>
<GID>679</GID>
<name>write_clock</name></connection>
<intersection>-212 9</intersection>
<intersection>-167.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-167.5,27,-167.5,82.5</points>
<intersection>27 7</intersection>
<intersection>82.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-212,27,-167.5,27</points>
<intersection>-212 8</intersection>
<intersection>-167.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-212,27,-212,40</points>
<connection>
<GID>460</GID>
<name>clock</name></connection>
<intersection>27 7</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-212,82.5,-212,87</points>
<intersection>82.5 1</intersection>
<intersection>87 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-212,87,-209,87</points>
<connection>
<GID>678</GID>
<name>IN_0</name></connection>
<intersection>-212 9</intersection></hsegment></shape></wire>
<wire>
<ID>573</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-224,81.5,-224,90</points>
<intersection>81.5 6</intersection>
<intersection>83.5 4</intersection>
<intersection>84.5 1</intersection>
<intersection>90 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-224,84.5,-222,84.5</points>
<connection>
<GID>679</GID>
<name>ADDRESS_7</name></connection>
<intersection>-224 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-232.5,90,-224,90</points>
<intersection>-232.5 9</intersection>
<intersection>-224 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-224,83.5,-222,83.5</points>
<connection>
<GID>679</GID>
<name>ADDRESS_6</name></connection>
<intersection>-224 0</intersection>
<intersection>-222 7</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-224,81.5,-222,81.5</points>
<connection>
<GID>679</GID>
<name>ADDRESS_4</name></connection>
<intersection>-224 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-222,82.5,-222,83.5</points>
<connection>
<GID>679</GID>
<name>ADDRESS_5</name></connection>
<intersection>83.5 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-232.5,89,-232.5,90</points>
<connection>
<GID>482</GID>
<name>OUT_0</name></connection>
<intersection>90 2</intersection></vsegment></shape></wire>
<wire>
<ID>577</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-212,79.5,-200,79.5</points>
<connection>
<GID>486</GID>
<name>OUT_0</name></connection>
<intersection>-212 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-212,79.5,-212,80.5</points>
<connection>
<GID>679</GID>
<name>ENABLE_0</name></connection>
<intersection>79.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>578</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-187,58,-187,64</points>
<connection>
<GID>638</GID>
<name>T_in2</name></connection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-198,58,-187,58</points>
<intersection>-198 2</intersection>
<intersection>-187 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-198,31,-198,58</points>
<intersection>31 3</intersection>
<intersection>42 6</intersection>
<intersection>58 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-198,31,-184.5,31</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<intersection>-198 2</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-207,42,-198,42</points>
<connection>
<GID>460</GID>
<name>OUT_0</name></connection>
<intersection>-198 2</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>6.575,-32.1253,161.375,-110.375</PageViewport>
<gate>
<ID>775</ID>
<type>AE_REGISTER8</type>
<position>31.5,-48.5</position>
<input>
<ID>IN_0</ID>713 </input>
<input>
<ID>IN_1</ID>714 </input>
<input>
<ID>IN_2</ID>715 </input>
<input>
<ID>IN_3</ID>716 </input>
<input>
<ID>IN_4</ID>717 </input>
<input>
<ID>IN_5</ID>718 </input>
<input>
<ID>IN_6</ID>719 </input>
<input>
<ID>IN_7</ID>720 </input>
<output>
<ID>OUT_0</ID>662 </output>
<output>
<ID>OUT_1</ID>657 </output>
<output>
<ID>OUT_2</ID>666 </output>
<output>
<ID>OUT_3</ID>694 </output>
<output>
<ID>OUT_4</ID>696 </output>
<output>
<ID>OUT_5</ID>699 </output>
<output>
<ID>OUT_6</ID>701 </output>
<output>
<ID>OUT_7</ID>705 </output>
<input>
<ID>clock</ID>712 </input>
<input>
<ID>load</ID>738 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>777</ID>
<type>AI_XOR2</type>
<position>42.5,-84.5</position>
<input>
<ID>IN_0</ID>662 </input>
<input>
<ID>IN_1</ID>581 </input>
<output>
<ID>OUT</ID>591 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>789</ID>
<type>AA_AND2</type>
<position>47.5,-79.5</position>
<input>
<ID>IN_0</ID>662 </input>
<input>
<ID>IN_1</ID>581 </input>
<output>
<ID>OUT</ID>648 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>799</ID>
<type>AI_XOR2</type>
<position>54.5,-78</position>
<input>
<ID>IN_0</ID>613 </input>
<input>
<ID>IN_1</ID>648 </input>
<output>
<ID>OUT</ID>649 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>801</ID>
<type>AA_AND2</type>
<position>54.5,-73</position>
<input>
<ID>IN_0</ID>613 </input>
<input>
<ID>IN_1</ID>648 </input>
<output>
<ID>OUT</ID>651 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>811</ID>
<type>AI_XOR2</type>
<position>54.5,-67</position>
<input>
<ID>IN_0</ID>657 </input>
<input>
<ID>IN_1</ID>649 </input>
<output>
<ID>OUT</ID>612 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>815</ID>
<type>AA_AND2</type>
<position>54.5,-62</position>
<input>
<ID>IN_0</ID>657 </input>
<input>
<ID>IN_1</ID>649 </input>
<output>
<ID>OUT</ID>650 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>817</ID>
<type>AE_REGISTER8</type>
<position>31,-95.5</position>
<input>
<ID>IN_0</ID>721 </input>
<input>
<ID>IN_1</ID>722 </input>
<input>
<ID>IN_2</ID>723 </input>
<input>
<ID>IN_3</ID>724 </input>
<input>
<ID>IN_4</ID>725 </input>
<input>
<ID>IN_5</ID>726 </input>
<input>
<ID>IN_6</ID>727 </input>
<input>
<ID>IN_7</ID>728 </input>
<output>
<ID>OUT_0</ID>581 </output>
<output>
<ID>OUT_1</ID>613 </output>
<output>
<ID>OUT_2</ID>614 </output>
<output>
<ID>OUT_3</ID>615 </output>
<output>
<ID>OUT_4</ID>616 </output>
<output>
<ID>OUT_5</ID>711 </output>
<output>
<ID>OUT_6</ID>640 </output>
<output>
<ID>OUT_7</ID>647 </output>
<input>
<ID>clock</ID>712 </input>
<input>
<ID>load</ID>739 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>819</ID>
<type>AE_REGISTER8</type>
<position>143.5,-87.5</position>
<input>
<ID>IN_0</ID>591 </input>
<input>
<ID>IN_1</ID>612 </input>
<input>
<ID>IN_2</ID>611 </input>
<input>
<ID>IN_3</ID>610 </input>
<input>
<ID>IN_4</ID>595 </input>
<input>
<ID>IN_5</ID>594 </input>
<input>
<ID>IN_6</ID>593 </input>
<input>
<ID>IN_7</ID>592 </input>
<output>
<ID>OUT_0</ID>736 </output>
<output>
<ID>OUT_1</ID>735 </output>
<output>
<ID>OUT_2</ID>734 </output>
<output>
<ID>OUT_3</ID>733 </output>
<output>
<ID>OUT_4</ID>732 </output>
<output>
<ID>OUT_5</ID>731 </output>
<output>
<ID>OUT_6</ID>730 </output>
<output>
<ID>OUT_7</ID>729 </output>
<input>
<ID>clock</ID>712 </input>
<input>
<ID>load</ID>740 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>820</ID>
<type>AE_OR2</type>
<position>54.5,-55</position>
<input>
<ID>IN_0</ID>651 </input>
<input>
<ID>IN_1</ID>650 </input>
<output>
<ID>OUT</ID>652 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>822</ID>
<type>AI_XOR2</type>
<position>68.5,-79.5</position>
<input>
<ID>IN_0</ID>652 </input>
<input>
<ID>IN_1</ID>614 </input>
<output>
<ID>OUT</ID>655 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>824</ID>
<type>AA_AND2</type>
<position>68.5,-74.5</position>
<input>
<ID>IN_0</ID>652 </input>
<input>
<ID>IN_1</ID>614 </input>
<output>
<ID>OUT</ID>654 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>825</ID>
<type>AI_XOR2</type>
<position>68.5,-68.5</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>655 </input>
<output>
<ID>OUT</ID>611 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>828</ID>
<type>AA_AND2</type>
<position>68.5,-63.5</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>655 </input>
<output>
<ID>OUT</ID>653 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>831</ID>
<type>AE_OR2</type>
<position>68.5,-56.5</position>
<input>
<ID>IN_0</ID>654 </input>
<input>
<ID>IN_1</ID>653 </input>
<output>
<ID>OUT</ID>656 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>860</ID>
<type>AI_XOR2</type>
<position>81.5,-79.5</position>
<input>
<ID>IN_0</ID>656 </input>
<input>
<ID>IN_1</ID>615 </input>
<output>
<ID>OUT</ID>661 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>861</ID>
<type>AA_AND2</type>
<position>81.5,-74.5</position>
<input>
<ID>IN_0</ID>656 </input>
<input>
<ID>IN_1</ID>615 </input>
<output>
<ID>OUT</ID>660 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>862</ID>
<type>AI_XOR2</type>
<position>81.5,-68.5</position>
<input>
<ID>IN_0</ID>694 </input>
<input>
<ID>IN_1</ID>661 </input>
<output>
<ID>OUT</ID>610 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>863</ID>
<type>AA_AND2</type>
<position>81.5,-63.5</position>
<input>
<ID>IN_0</ID>694 </input>
<input>
<ID>IN_1</ID>661 </input>
<output>
<ID>OUT</ID>659 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>864</ID>
<type>AE_OR2</type>
<position>81.5,-56.5</position>
<input>
<ID>IN_0</ID>660 </input>
<input>
<ID>IN_1</ID>659 </input>
<output>
<ID>OUT</ID>664 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>865</ID>
<type>AI_XOR2</type>
<position>94,-79.5</position>
<input>
<ID>IN_0</ID>664 </input>
<input>
<ID>IN_1</ID>616 </input>
<output>
<ID>OUT</ID>737 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>866</ID>
<type>AA_AND2</type>
<position>94,-74.5</position>
<input>
<ID>IN_0</ID>664 </input>
<input>
<ID>IN_1</ID>616 </input>
<output>
<ID>OUT</ID>693 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>867</ID>
<type>AI_XOR2</type>
<position>94,-68.5</position>
<input>
<ID>IN_0</ID>696 </input>
<input>
<ID>IN_1</ID>737 </input>
<output>
<ID>OUT</ID>595 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>868</ID>
<type>AA_AND2</type>
<position>94,-63.5</position>
<input>
<ID>IN_0</ID>696 </input>
<input>
<ID>IN_1</ID>737 </input>
<output>
<ID>OUT</ID>692 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>869</ID>
<type>AE_OR2</type>
<position>94,-56.5</position>
<input>
<ID>IN_0</ID>693 </input>
<input>
<ID>IN_1</ID>692 </input>
<output>
<ID>OUT</ID>695 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>870</ID>
<type>AI_XOR2</type>
<position>107,-79.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>711 </input>
<output>
<ID>OUT</ID>709 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>872</ID>
<type>AA_AND2</type>
<position>107,-74.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>711 </input>
<output>
<ID>OUT</ID>698 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>873</ID>
<type>AI_XOR2</type>
<position>107,-68.5</position>
<input>
<ID>IN_0</ID>699 </input>
<input>
<ID>IN_1</ID>709 </input>
<output>
<ID>OUT</ID>594 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>874</ID>
<type>AA_AND2</type>
<position>107,-63.5</position>
<input>
<ID>IN_0</ID>699 </input>
<input>
<ID>IN_1</ID>709 </input>
<output>
<ID>OUT</ID>697 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>875</ID>
<type>AE_OR2</type>
<position>107,-56.5</position>
<input>
<ID>IN_0</ID>698 </input>
<input>
<ID>IN_1</ID>697 </input>
<output>
<ID>OUT</ID>700 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>876</ID>
<type>AI_XOR2</type>
<position>120,-79.5</position>
<input>
<ID>IN_0</ID>700 </input>
<input>
<ID>IN_1</ID>640 </input>
<output>
<ID>OUT</ID>704 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>877</ID>
<type>AA_AND2</type>
<position>120,-74.5</position>
<input>
<ID>IN_0</ID>700 </input>
<input>
<ID>IN_1</ID>640 </input>
<output>
<ID>OUT</ID>703 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>878</ID>
<type>AI_XOR2</type>
<position>120,-68.5</position>
<input>
<ID>IN_0</ID>701 </input>
<input>
<ID>IN_1</ID>704 </input>
<output>
<ID>OUT</ID>593 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>879</ID>
<type>AA_AND2</type>
<position>120,-63.5</position>
<input>
<ID>IN_0</ID>701 </input>
<input>
<ID>IN_1</ID>704 </input>
<output>
<ID>OUT</ID>702 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>880</ID>
<type>AE_OR2</type>
<position>120,-56.5</position>
<input>
<ID>IN_0</ID>703 </input>
<input>
<ID>IN_1</ID>702 </input>
<output>
<ID>OUT</ID>706 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>881</ID>
<type>AI_XOR2</type>
<position>132.5,-79.5</position>
<input>
<ID>IN_0</ID>706 </input>
<input>
<ID>IN_1</ID>647 </input>
<output>
<ID>OUT</ID>710 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>882</ID>
<type>AA_AND2</type>
<position>132.5,-74.5</position>
<input>
<ID>IN_0</ID>706 </input>
<input>
<ID>IN_1</ID>647 </input>
<output>
<ID>OUT</ID>708 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>883</ID>
<type>AI_XOR2</type>
<position>132.5,-68.5</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>710 </input>
<output>
<ID>OUT</ID>592 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>691</ID>
<type>DA_FROM</type>
<position>26.5,-36</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-ADDER</lparam></gate>
<gate>
<ID>884</ID>
<type>AA_AND2</type>
<position>132.5,-63.5</position>
<input>
<ID>IN_0</ID>705 </input>
<input>
<ID>IN_1</ID>710 </input>
<output>
<ID>OUT</ID>707 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>692</ID>
<type>DA_FROM</type>
<position>26.5,-83.5</position>
<input>
<ID>IN_0</ID>739 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-ADDER</lparam></gate>
<gate>
<ID>885</ID>
<type>AE_OR2</type>
<position>132.5,-56.5</position>
<input>
<ID>IN_0</ID>708 </input>
<input>
<ID>IN_1</ID>707 </input>
<output>
<ID>OUT</ID>617 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>693</ID>
<type>DA_FROM</type>
<position>159,-73</position>
<input>
<ID>IN_0</ID>740 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID LOAD-ADDER-RESULT</lparam></gate>
<gate>
<ID>886</ID>
<type>AA_LABEL</type>
<position>85.5,-37</position>
<gparam>LABEL_TEXT 8-bit Adder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>694</ID>
<type>DA_FROM</type>
<position>36.5,-106.5</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK-PULSE-IN</lparam></gate>
<gate>
<ID>695</ID>
<type>DE_TO</type>
<position>137.5,-56.5</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-OVERFLOW</lparam></gate>
<gate>
<ID>696</ID>
<type>DA_FROM</type>
<position>19.5,-40</position>
<input>
<ID>IN_0</ID>720 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-7</lparam></gate>
<gate>
<ID>697</ID>
<type>DA_FROM</type>
<position>19.5,-42</position>
<input>
<ID>IN_0</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-6</lparam></gate>
<gate>
<ID>698</ID>
<type>DA_FROM</type>
<position>19.5,-44</position>
<input>
<ID>IN_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-5</lparam></gate>
<gate>
<ID>699</ID>
<type>DA_FROM</type>
<position>19.5,-46</position>
<input>
<ID>IN_0</ID>717 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-4</lparam></gate>
<gate>
<ID>700</ID>
<type>DA_FROM</type>
<position>19.5,-48</position>
<input>
<ID>IN_0</ID>716 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-3</lparam></gate>
<gate>
<ID>701</ID>
<type>DA_FROM</type>
<position>19.5,-50</position>
<input>
<ID>IN_0</ID>715 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-2</lparam></gate>
<gate>
<ID>702</ID>
<type>DA_FROM</type>
<position>19.5,-52</position>
<input>
<ID>IN_0</ID>714 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-1</lparam></gate>
<gate>
<ID>703</ID>
<type>DA_FROM</type>
<position>19.5,-54</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-0</lparam></gate>
<gate>
<ID>704</ID>
<type>DA_FROM</type>
<position>19.5,-87.5</position>
<input>
<ID>IN_0</ID>728 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-7</lparam></gate>
<gate>
<ID>705</ID>
<type>DA_FROM</type>
<position>19.5,-89.5</position>
<input>
<ID>IN_0</ID>727 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-6</lparam></gate>
<gate>
<ID>706</ID>
<type>DA_FROM</type>
<position>19.5,-91.5</position>
<input>
<ID>IN_0</ID>726 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-5</lparam></gate>
<gate>
<ID>707</ID>
<type>DA_FROM</type>
<position>19.5,-93.5</position>
<input>
<ID>IN_0</ID>725 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-4</lparam></gate>
<gate>
<ID>708</ID>
<type>DA_FROM</type>
<position>19.5,-95.5</position>
<input>
<ID>IN_0</ID>724 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-3</lparam></gate>
<gate>
<ID>710</ID>
<type>DA_FROM</type>
<position>19.5,-97.5</position>
<input>
<ID>IN_0</ID>723 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-2</lparam></gate>
<gate>
<ID>713</ID>
<type>DA_FROM</type>
<position>19.5,-99.5</position>
<input>
<ID>IN_0</ID>722 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-1</lparam></gate>
<gate>
<ID>725</ID>
<type>DA_FROM</type>
<position>19.5,-101.5</position>
<input>
<ID>IN_0</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-0</lparam></gate>
<gate>
<ID>729</ID>
<type>DE_TO</type>
<position>154,-80</position>
<input>
<ID>IN_0</ID>729 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-7</lparam></gate>
<gate>
<ID>759</ID>
<type>DE_TO</type>
<position>154,-82</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-6</lparam></gate>
<gate>
<ID>762</ID>
<type>DE_TO</type>
<position>154,-84</position>
<input>
<ID>IN_0</ID>731 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-5</lparam></gate>
<gate>
<ID>765</ID>
<type>DE_TO</type>
<position>154,-86</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-4</lparam></gate>
<gate>
<ID>766</ID>
<type>DE_TO</type>
<position>154,-88</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-3</lparam></gate>
<gate>
<ID>767</ID>
<type>DE_TO</type>
<position>154,-90</position>
<input>
<ID>IN_0</ID>734 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-2</lparam></gate>
<gate>
<ID>768</ID>
<type>DE_TO</type>
<position>154,-92</position>
<input>
<ID>IN_0</ID>735 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-1</lparam></gate>
<gate>
<ID>770</ID>
<type>DE_TO</type>
<position>154,-94</position>
<input>
<ID>IN_0</ID>736 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-0</lparam></gate>
<wire>
<ID>581</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-98.5,38.5,-80.5</points>
<intersection>-98.5 4</intersection>
<intersection>-85.5 2</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-80.5,44.5,-80.5</points>
<connection>
<GID>789</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-85.5,39.5,-85.5</points>
<connection>
<GID>777</GID>
<name>IN_1</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35,-98.5,38.5,-98.5</points>
<connection>
<GID>817</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>591</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-90.5,46.5,-84.5</points>
<intersection>-90.5 2</intersection>
<intersection>-84.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-84.5,46.5,-84.5</points>
<connection>
<GID>777</GID>
<name>OUT</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-90.5,139.5,-90.5</points>
<connection>
<GID>819</GID>
<name>IN_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>592</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,-83.5,137,-68.5</points>
<intersection>-83.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-68.5,137,-68.5</points>
<connection>
<GID>883</GID>
<name>OUT</name></connection>
<intersection>137 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137,-83.5,139.5,-83.5</points>
<connection>
<GID>819</GID>
<name>IN_7</name></connection>
<intersection>137 0</intersection></hsegment></shape></wire>
<wire>
<ID>593</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-84.5,124.5,-68.5</points>
<intersection>-84.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-68.5,124.5,-68.5</points>
<connection>
<GID>878</GID>
<name>OUT</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-84.5,139.5,-84.5</points>
<connection>
<GID>819</GID>
<name>IN_6</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>594</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-85.5,110.5,-68.5</points>
<intersection>-85.5 6</intersection>
<intersection>-68.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>110,-68.5,110.5,-68.5</points>
<connection>
<GID>873</GID>
<name>OUT</name></connection>
<intersection>110.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>110.5,-85.5,139.5,-85.5</points>
<connection>
<GID>819</GID>
<name>IN_5</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>595</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-86.5,97.5,-68.5</points>
<intersection>-86.5 5</intersection>
<intersection>-68.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>97,-68.5,97.5,-68.5</points>
<connection>
<GID>867</GID>
<name>OUT</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>97.5,-86.5,139.5,-86.5</points>
<connection>
<GID>819</GID>
<name>IN_4</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>610</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-87.5,84.5,-68.5</points>
<connection>
<GID>862</GID>
<name>OUT</name></connection>
<intersection>-87.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>84.5,-87.5,139.5,-87.5</points>
<connection>
<GID>819</GID>
<name>IN_3</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>611</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-88.5,72,-68.5</points>
<intersection>-88.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-68.5,72,-68.5</points>
<connection>
<GID>825</GID>
<name>OUT</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-88.5,139.5,-88.5</points>
<connection>
<GID>819</GID>
<name>IN_2</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>612</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-89.5,60.5,-67</points>
<intersection>-89.5 4</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57.5,-67,60.5,-67</points>
<connection>
<GID>811</GID>
<name>OUT</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>60.5,-89.5,139.5,-89.5</points>
<connection>
<GID>819</GID>
<name>IN_1</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>613</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-97.5,37.5,-72</points>
<intersection>-97.5 3</intersection>
<intersection>-77 5</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-72,51.5,-72</points>
<connection>
<GID>801</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>35,-97.5,37.5,-97.5</points>
<connection>
<GID>817</GID>
<name>OUT_1</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>37.5,-77,51.5,-77</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>614</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-96.5,61.5,-75.5</points>
<intersection>-96.5 1</intersection>
<intersection>-80.5 3</intersection>
<intersection>-75.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-96.5,61.5,-96.5</points>
<connection>
<GID>817</GID>
<name>OUT_2</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-75.5,65.5,-75.5</points>
<connection>
<GID>824</GID>
<name>IN_1</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>61.5,-80.5,65.5,-80.5</points>
<connection>
<GID>822</GID>
<name>IN_1</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>615</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-95.5,74.5,-80.5</points>
<intersection>-95.5 2</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-80.5,78.5,-80.5</points>
<connection>
<GID>860</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection>
<intersection>77 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-95.5,74.5,-95.5</points>
<connection>
<GID>817</GID>
<name>OUT_3</name></connection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77,-80.5,77,-75.5</points>
<intersection>-80.5 1</intersection>
<intersection>-75.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>77,-75.5,78.5,-75.5</points>
<connection>
<GID>861</GID>
<name>IN_1</name></connection>
<intersection>77 3</intersection></hsegment></shape></wire>
<wire>
<ID>616</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-94.5,85.5,-80.5</points>
<intersection>-94.5 12</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-80.5,91,-80.5</points>
<connection>
<GID>865</GID>
<name>IN_1</name></connection>
<intersection>85.5 0</intersection>
<intersection>89.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89.5,-80.5,89.5,-75.5</points>
<intersection>-80.5 1</intersection>
<intersection>-75.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>89.5,-75.5,91,-75.5</points>
<connection>
<GID>866</GID>
<name>IN_1</name></connection>
<intersection>89.5 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>35,-94.5,85.5,-94.5</points>
<connection>
<GID>817</GID>
<name>OUT_4</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>617</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-56.5,135.5,-56.5</points>
<connection>
<GID>885</GID>
<name>OUT</name></connection>
<connection>
<GID>695</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>640</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109.5,-92.5,109.5,-80.5</points>
<intersection>-92.5 7</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>109.5,-80.5,117,-80.5</points>
<connection>
<GID>876</GID>
<name>IN_1</name></connection>
<intersection>109.5 0</intersection>
<intersection>115.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-80.5,115.5,-75.5</points>
<intersection>-80.5 1</intersection>
<intersection>-75.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>115.5,-75.5,117,-75.5</points>
<connection>
<GID>877</GID>
<name>IN_1</name></connection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>35,-92.5,109.5,-92.5</points>
<connection>
<GID>817</GID>
<name>OUT_6</name></connection>
<intersection>109.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>647</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-91.5,123,-80.5</points>
<intersection>-91.5 5</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-80.5,129.5,-80.5</points>
<connection>
<GID>881</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection>
<intersection>128.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,-80.5,128.5,-75.5</points>
<intersection>-80.5 1</intersection>
<intersection>-75.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>128.5,-75.5,129.5,-75.5</points>
<connection>
<GID>882</GID>
<name>IN_1</name></connection>
<intersection>128.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>35,-91.5,123,-91.5</points>
<connection>
<GID>817</GID>
<name>OUT_7</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>648</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-79.5,50.5,-74</points>
<connection>
<GID>789</GID>
<name>OUT</name></connection>
<intersection>-79 1</intersection>
<intersection>-74 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-79,51.5,-79</points>
<connection>
<GID>799</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-74,51.5,-74</points>
<connection>
<GID>801</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>649</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-78,59.5,-69.5</points>
<intersection>-78 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-69.5,59.5,-69.5</points>
<intersection>51 3</intersection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-78,59.5,-78</points>
<connection>
<GID>799</GID>
<name>OUT</name></connection>
<intersection>59.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51,-69.5,51,-63</points>
<intersection>-69.5 1</intersection>
<intersection>-68 4</intersection>
<intersection>-63 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>51,-68,51.5,-68</points>
<connection>
<GID>811</GID>
<name>IN_1</name></connection>
<intersection>51 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>51,-63,51.5,-63</points>
<connection>
<GID>815</GID>
<name>IN_1</name></connection>
<intersection>51 3</intersection></hsegment></shape></wire>
<wire>
<ID>650</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>51.5,-59.5,57.5,-59.5</points>
<intersection>51.5 4</intersection>
<intersection>57.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57.5,-62,57.5,-59.5</points>
<connection>
<GID>815</GID>
<name>OUT</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>51.5,-59.5,51.5,-56</points>
<connection>
<GID>820</GID>
<name>IN_1</name></connection>
<intersection>-59.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>651</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-58,58.5,-58</points>
<intersection>49.5 4</intersection>
<intersection>58.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58.5,-73,58.5,-58</points>
<intersection>-73 6</intersection>
<intersection>-58 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>49.5,-58,49.5,-54</points>
<intersection>-58 1</intersection>
<intersection>-54 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>49.5,-54,51.5,-54</points>
<connection>
<GID>820</GID>
<name>IN_0</name></connection>
<intersection>49.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>57.5,-73,58.5,-73</points>
<connection>
<GID>801</GID>
<name>OUT</name></connection>
<intersection>58.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>652</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>62,-78.5,62,-55</points>
<intersection>-78.5 8</intersection>
<intersection>-73.5 9</intersection>
<intersection>-55 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>57.5,-55,62,-55</points>
<connection>
<GID>820</GID>
<name>OUT</name></connection>
<intersection>62 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>62,-78.5,65.5,-78.5</points>
<connection>
<GID>822</GID>
<name>IN_0</name></connection>
<intersection>62 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>62,-73.5,65.5,-73.5</points>
<connection>
<GID>824</GID>
<name>IN_0</name></connection>
<intersection>62 5</intersection></hsegment></shape></wire>
<wire>
<ID>653</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>65.5,-61,71.5,-61</points>
<intersection>65.5 4</intersection>
<intersection>71.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71.5,-63.5,71.5,-61</points>
<connection>
<GID>828</GID>
<name>OUT</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>65.5,-61,65.5,-57.5</points>
<connection>
<GID>831</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment></shape></wire>
<wire>
<ID>654</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63.5,-59.5,72.5,-59.5</points>
<intersection>63.5 4</intersection>
<intersection>72.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72.5,-74.5,72.5,-59.5</points>
<intersection>-74.5 6</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>63.5,-59.5,63.5,-55.5</points>
<intersection>-59.5 1</intersection>
<intersection>-55.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>63.5,-55.5,65.5,-55.5</points>
<connection>
<GID>831</GID>
<name>IN_0</name></connection>
<intersection>63.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>71.5,-74.5,72.5,-74.5</points>
<connection>
<GID>824</GID>
<name>OUT</name></connection>
<intersection>72.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>655</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-79.5,73.5,-71.5</points>
<intersection>-79.5 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-71.5,73.5,-71.5</points>
<intersection>64 3</intersection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,-79.5,73.5,-79.5</points>
<connection>
<GID>822</GID>
<name>OUT</name></connection>
<intersection>73.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>64,-71.5,64,-64.5</points>
<intersection>-71.5 1</intersection>
<intersection>-69.5 12</intersection>
<intersection>-64.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>64,-64.5,65.5,-64.5</points>
<connection>
<GID>828</GID>
<name>IN_1</name></connection>
<intersection>64 3</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>64,-69.5,65.5,-69.5</points>
<connection>
<GID>825</GID>
<name>IN_1</name></connection>
<intersection>64 3</intersection></hsegment></shape></wire>
<wire>
<ID>656</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>75,-78.5,75,-56.5</points>
<intersection>-78.5 8</intersection>
<intersection>-73.5 9</intersection>
<intersection>-56.5 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>75,-78.5,78.5,-78.5</points>
<connection>
<GID>860</GID>
<name>IN_0</name></connection>
<intersection>75 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>75,-73.5,78.5,-73.5</points>
<connection>
<GID>861</GID>
<name>IN_0</name></connection>
<intersection>75 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>71.5,-56.5,75,-56.5</points>
<connection>
<GID>831</GID>
<name>OUT</name></connection>
<intersection>75 5</intersection></hsegment></shape></wire>
<wire>
<ID>657</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>47.5,-66,47.5,-50.5</points>
<intersection>-66 6</intersection>
<intersection>-61 4</intersection>
<intersection>-50.5 7</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47.5,-61,51.5,-61</points>
<connection>
<GID>815</GID>
<name>IN_0</name></connection>
<intersection>47.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>47.5,-66,51.5,-66</points>
<connection>
<GID>811</GID>
<name>IN_0</name></connection>
<intersection>47.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>35.5,-50.5,47.5,-50.5</points>
<connection>
<GID>775</GID>
<name>OUT_1</name></connection>
<intersection>47.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>659</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-61,84.5,-61</points>
<intersection>78 4</intersection>
<intersection>84.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84.5,-63.5,84.5,-61</points>
<connection>
<GID>863</GID>
<name>OUT</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>78,-61,78,-57.5</points>
<intersection>-61 1</intersection>
<intersection>-57.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>78,-57.5,78.5,-57.5</points>
<connection>
<GID>864</GID>
<name>IN_1</name></connection>
<intersection>78 4</intersection></hsegment></shape></wire>
<wire>
<ID>660</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,-59.5,86,-59.5</points>
<intersection>77 4</intersection>
<intersection>86 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>86,-74.5,86,-59.5</points>
<intersection>-74.5 6</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>77,-59.5,77,-55.5</points>
<intersection>-59.5 1</intersection>
<intersection>-55.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>77,-55.5,78.5,-55.5</points>
<connection>
<GID>864</GID>
<name>IN_0</name></connection>
<intersection>77 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>84.5,-74.5,86,-74.5</points>
<connection>
<GID>861</GID>
<name>OUT</name></connection>
<intersection>86 3</intersection></hsegment></shape></wire>
<wire>
<ID>661</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-79.5,86.5,-71.5</points>
<intersection>-79.5 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-71.5,86.5,-71.5</points>
<intersection>77 3</intersection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-79.5,86.5,-79.5</points>
<connection>
<GID>860</GID>
<name>OUT</name></connection>
<intersection>86.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>77,-71.5,77,-64.5</points>
<intersection>-71.5 1</intersection>
<intersection>-69.5 9</intersection>
<intersection>-64.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>77,-64.5,78.5,-64.5</points>
<connection>
<GID>863</GID>
<name>IN_1</name></connection>
<intersection>77 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>77,-69.5,78.5,-69.5</points>
<connection>
<GID>862</GID>
<name>IN_1</name></connection>
<intersection>77 3</intersection></hsegment></shape></wire>
<wire>
<ID>662</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>35.5,-83.5,35.5,-51.5</points>
<connection>
<GID>775</GID>
<name>OUT_0</name></connection>
<intersection>-83.5 7</intersection>
<intersection>-78.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>35.5,-78.5,44.5,-78.5</points>
<connection>
<GID>789</GID>
<name>IN_0</name></connection>
<intersection>35.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>35.5,-83.5,39.5,-83.5</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<intersection>35.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>664</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>87.5,-78.5,87.5,-56.5</points>
<intersection>-78.5 8</intersection>
<intersection>-73.5 9</intersection>
<intersection>-56.5 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>87.5,-78.5,91,-78.5</points>
<connection>
<GID>865</GID>
<name>IN_0</name></connection>
<intersection>87.5 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>87.5,-73.5,91,-73.5</points>
<connection>
<GID>866</GID>
<name>IN_0</name></connection>
<intersection>87.5 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>84.5,-56.5,87.5,-56.5</points>
<connection>
<GID>864</GID>
<name>OUT</name></connection>
<intersection>87.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>666</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-67.5,63,-49.5</points>
<intersection>-67.5 2</intersection>
<intersection>-62.5 3</intersection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-49.5,63,-49.5</points>
<connection>
<GID>775</GID>
<name>OUT_2</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-67.5,65.5,-67.5</points>
<connection>
<GID>825</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>63,-62.5,65.5,-62.5</points>
<connection>
<GID>828</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>692</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-61,97,-61</points>
<intersection>90.5 4</intersection>
<intersection>97 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97,-63.5,97,-61</points>
<connection>
<GID>868</GID>
<name>OUT</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>90.5,-61,90.5,-57.5</points>
<intersection>-61 1</intersection>
<intersection>-57.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>90.5,-57.5,91,-57.5</points>
<connection>
<GID>869</GID>
<name>IN_1</name></connection>
<intersection>90.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>693</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-59.5,98.5,-59.5</points>
<intersection>89.5 4</intersection>
<intersection>98.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>98.5,-74.5,98.5,-59.5</points>
<intersection>-74.5 6</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>89.5,-59.5,89.5,-55.5</points>
<intersection>-59.5 1</intersection>
<intersection>-55.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>89.5,-55.5,91,-55.5</points>
<connection>
<GID>869</GID>
<name>IN_0</name></connection>
<intersection>89.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>97,-74.5,98.5,-74.5</points>
<connection>
<GID>866</GID>
<name>OUT</name></connection>
<intersection>98.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>694</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-67.5,76,-48.5</points>
<intersection>-67.5 2</intersection>
<intersection>-62.5 3</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-48.5,76,-48.5</points>
<connection>
<GID>775</GID>
<name>OUT_3</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-67.5,78.5,-67.5</points>
<connection>
<GID>862</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>76,-62.5,78.5,-62.5</points>
<connection>
<GID>863</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>695</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>100,-78.5,100,-56.5</points>
<intersection>-78.5 8</intersection>
<intersection>-73.5 9</intersection>
<intersection>-56.5 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>100,-78.5,104,-78.5</points>
<connection>
<GID>870</GID>
<name>IN_0</name></connection>
<intersection>100 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>100,-73.5,104,-73.5</points>
<connection>
<GID>872</GID>
<name>IN_0</name></connection>
<intersection>100 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>97,-56.5,100,-56.5</points>
<connection>
<GID>869</GID>
<name>OUT</name></connection>
<intersection>100 5</intersection></hsegment></shape></wire>
<wire>
<ID>696</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-67.5,88.5,-47.5</points>
<intersection>-67.5 2</intersection>
<intersection>-62.5 3</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-47.5,88.5,-47.5</points>
<connection>
<GID>775</GID>
<name>OUT_4</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88.5,-67.5,91,-67.5</points>
<connection>
<GID>867</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>88.5,-62.5,91,-62.5</points>
<connection>
<GID>868</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>697</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-61,110,-61</points>
<intersection>104 4</intersection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,-63.5,110,-61</points>
<connection>
<GID>874</GID>
<name>OUT</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>104,-61,104,-57.5</points>
<connection>
<GID>875</GID>
<name>IN_1</name></connection>
<intersection>-61 1</intersection></vsegment></shape></wire>
<wire>
<ID>698</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>102,-59.5,111,-59.5</points>
<intersection>102 4</intersection>
<intersection>111 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,-74.5,111,-59.5</points>
<intersection>-74.5 6</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>102,-59.5,102,-55.5</points>
<intersection>-59.5 1</intersection>
<intersection>-55.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>102,-55.5,104,-55.5</points>
<connection>
<GID>875</GID>
<name>IN_0</name></connection>
<intersection>102 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>110,-74.5,111,-74.5</points>
<connection>
<GID>872</GID>
<name>OUT</name></connection>
<intersection>111 3</intersection></hsegment></shape></wire>
<wire>
<ID>699</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-67.5,101.5,-46.5</points>
<intersection>-67.5 2</intersection>
<intersection>-62.5 3</intersection>
<intersection>-46.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>101.5,-67.5,104,-67.5</points>
<connection>
<GID>873</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>101.5,-62.5,104,-62.5</points>
<connection>
<GID>874</GID>
<name>IN_0</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35.5,-46.5,101.5,-46.5</points>
<connection>
<GID>775</GID>
<name>OUT_5</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>700</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>113.5,-78.5,113.5,-56.5</points>
<intersection>-78.5 8</intersection>
<intersection>-73.5 9</intersection>
<intersection>-56.5 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>113.5,-78.5,117,-78.5</points>
<connection>
<GID>876</GID>
<name>IN_0</name></connection>
<intersection>113.5 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>113.5,-73.5,117,-73.5</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<intersection>113.5 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>110,-56.5,113.5,-56.5</points>
<connection>
<GID>875</GID>
<name>OUT</name></connection>
<intersection>113.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>701</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-67.5,114.5,-45.5</points>
<intersection>-67.5 2</intersection>
<intersection>-62.5 3</intersection>
<intersection>-45.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-67.5,117,-67.5</points>
<connection>
<GID>878</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>114.5,-62.5,117,-62.5</points>
<connection>
<GID>879</GID>
<name>IN_0</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35.5,-45.5,114.5,-45.5</points>
<connection>
<GID>775</GID>
<name>OUT_6</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>702</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,-61,123,-61</points>
<intersection>116.5 4</intersection>
<intersection>123 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>123,-63.5,123,-61</points>
<connection>
<GID>879</GID>
<name>OUT</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>116.5,-61,116.5,-57.5</points>
<intersection>-61 1</intersection>
<intersection>-57.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>116.5,-57.5,117,-57.5</points>
<connection>
<GID>880</GID>
<name>IN_1</name></connection>
<intersection>116.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>703</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115.5,-59.5,124.5,-59.5</points>
<intersection>115.5 4</intersection>
<intersection>124.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>124.5,-74.5,124.5,-59.5</points>
<intersection>-74.5 6</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>115.5,-59.5,115.5,-55.5</points>
<intersection>-59.5 1</intersection>
<intersection>-55.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>115.5,-55.5,117,-55.5</points>
<connection>
<GID>880</GID>
<name>IN_0</name></connection>
<intersection>115.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>123,-74.5,124.5,-74.5</points>
<connection>
<GID>877</GID>
<name>OUT</name></connection>
<intersection>124.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>704</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-79.5,125,-71.5</points>
<intersection>-79.5 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-71.5,125,-71.5</points>
<intersection>115.5 3</intersection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123,-79.5,125,-79.5</points>
<connection>
<GID>876</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115.5,-71.5,115.5,-64.5</points>
<intersection>-71.5 1</intersection>
<intersection>-69.5 9</intersection>
<intersection>-64.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>115.5,-64.5,117,-64.5</points>
<connection>
<GID>879</GID>
<name>IN_1</name></connection>
<intersection>115.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>115.5,-69.5,117,-69.5</points>
<connection>
<GID>878</GID>
<name>IN_1</name></connection>
<intersection>115.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>705</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-67.5,127,-44.5</points>
<intersection>-67.5 2</intersection>
<intersection>-62.5 3</intersection>
<intersection>-44.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>127,-67.5,129.5,-67.5</points>
<connection>
<GID>883</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>127,-62.5,129.5,-62.5</points>
<connection>
<GID>884</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35.5,-44.5,127,-44.5</points>
<connection>
<GID>775</GID>
<name>OUT_7</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>706</ID>
<shape>
<vsegment>
<ID>5</ID>
<points>126,-78.5,126,-56.5</points>
<intersection>-78.5 8</intersection>
<intersection>-73.5 9</intersection>
<intersection>-56.5 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>126,-78.5,129.5,-78.5</points>
<connection>
<GID>881</GID>
<name>IN_0</name></connection>
<intersection>126 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>126,-73.5,129.5,-73.5</points>
<connection>
<GID>882</GID>
<name>IN_0</name></connection>
<intersection>126 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>123,-56.5,126,-56.5</points>
<connection>
<GID>880</GID>
<name>OUT</name></connection>
<intersection>126 5</intersection></hsegment></shape></wire>
<wire>
<ID>707</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129,-61,135.5,-61</points>
<intersection>129 4</intersection>
<intersection>135.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>135.5,-63.5,135.5,-61</points>
<connection>
<GID>884</GID>
<name>OUT</name></connection>
<intersection>-61 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>129,-61,129,-57.5</points>
<intersection>-61 1</intersection>
<intersection>-57.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>129,-57.5,129.5,-57.5</points>
<connection>
<GID>885</GID>
<name>IN_1</name></connection>
<intersection>129 4</intersection></hsegment></shape></wire>
<wire>
<ID>708</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>128,-59.5,138,-59.5</points>
<intersection>128 4</intersection>
<intersection>138 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>138,-74.5,138,-59.5</points>
<intersection>-74.5 6</intersection>
<intersection>-59.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>128,-59.5,128,-55.5</points>
<intersection>-59.5 1</intersection>
<intersection>-55.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>128,-55.5,129.5,-55.5</points>
<connection>
<GID>885</GID>
<name>IN_0</name></connection>
<intersection>128 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>135.5,-74.5,138,-74.5</points>
<connection>
<GID>882</GID>
<name>OUT</name></connection>
<intersection>138 3</intersection></hsegment></shape></wire>
<wire>
<ID>709</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-79.5,112,-71.5</points>
<intersection>-79.5 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-71.5,112,-71.5</points>
<intersection>103 3</intersection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-79.5,112,-79.5</points>
<connection>
<GID>870</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103,-71.5,103,-64.5</points>
<intersection>-71.5 1</intersection>
<intersection>-69.5 6</intersection>
<intersection>-64.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>103,-64.5,104,-64.5</points>
<connection>
<GID>874</GID>
<name>IN_1</name></connection>
<intersection>103 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>103,-69.5,104,-69.5</points>
<connection>
<GID>873</GID>
<name>IN_1</name></connection>
<intersection>103 3</intersection></hsegment></shape></wire>
<wire>
<ID>710</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-79.5,136,-71.5</points>
<intersection>-79.5 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,-71.5,136,-71.5</points>
<intersection>128.5 3</intersection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>135.5,-79.5,136,-79.5</points>
<connection>
<GID>881</GID>
<name>OUT</name></connection>
<intersection>136 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,-71.5,128.5,-64.5</points>
<intersection>-71.5 1</intersection>
<intersection>-69.5 4</intersection>
<intersection>-64.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>128.5,-69.5,129.5,-69.5</points>
<connection>
<GID>883</GID>
<name>IN_1</name></connection>
<intersection>128.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>128.5,-64.5,129.5,-64.5</points>
<connection>
<GID>884</GID>
<name>IN_1</name></connection>
<intersection>128.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>711</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-93.5,99.5,-80.5</points>
<intersection>-93.5 2</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-80.5,104,-80.5</points>
<connection>
<GID>870</GID>
<name>IN_1</name></connection>
<intersection>99.5 0</intersection>
<intersection>102 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-93.5,99.5,-93.5</points>
<connection>
<GID>817</GID>
<name>OUT_5</name></connection>
<intersection>99.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>102,-80.5,102,-75.5</points>
<intersection>-80.5 1</intersection>
<intersection>-75.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>102,-75.5,104,-75.5</points>
<connection>
<GID>872</GID>
<name>IN_1</name></connection>
<intersection>102 3</intersection></hsegment></shape></wire>
<wire>
<ID>712</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-106.5,43,-56</points>
<intersection>-106.5 3</intersection>
<intersection>-103 6</intersection>
<intersection>-56 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>38.5,-106.5,142.5,-106.5</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection>
<intersection>142.5 5</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>30.5,-56,43,-56</points>
<intersection>30.5 8</intersection>
<intersection>43 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>142.5,-106.5,142.5,-92.5</points>
<connection>
<GID>819</GID>
<name>clock</name></connection>
<intersection>-106.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>30,-103,43,-103</points>
<intersection>30 7</intersection>
<intersection>43 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>30,-103,30,-100.5</points>
<connection>
<GID>817</GID>
<name>clock</name></connection>
<intersection>-103 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>30.5,-56,30.5,-53.5</points>
<connection>
<GID>775</GID>
<name>clock</name></connection>
<intersection>-56 4</intersection></vsegment></shape></wire>
<wire>
<ID>713</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-54,27.5,-51.5</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-54,27.5,-54</points>
<connection>
<GID>703</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>714</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-52,26.5,-50.5</points>
<intersection>-52 2</intersection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-50.5,27.5,-50.5</points>
<connection>
<GID>775</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-52,26.5,-52</points>
<connection>
<GID>702</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>715</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-50,24.5,-49.5</points>
<intersection>-50 2</intersection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-49.5,27.5,-49.5</points>
<connection>
<GID>775</GID>
<name>IN_2</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-50,24.5,-50</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>716</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-48.5,27.5,-48.5</points>
<connection>
<GID>775</GID>
<name>IN_3</name></connection>
<intersection>21.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-48.5,21.5,-48</points>
<connection>
<GID>700</GID>
<name>IN_0</name></connection>
<intersection>-48.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>717</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-47.5,22,-46</points>
<intersection>-47.5 1</intersection>
<intersection>-46 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-47.5,27.5,-47.5</points>
<connection>
<GID>775</GID>
<name>IN_4</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>21.5,-46,22,-46</points>
<connection>
<GID>699</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>718</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-46.5,22.5,-44</points>
<intersection>-46.5 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-46.5,27.5,-46.5</points>
<connection>
<GID>775</GID>
<name>IN_5</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-44,22.5,-44</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>719</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-45.5,23.5,-42</points>
<intersection>-45.5 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-45.5,27.5,-45.5</points>
<connection>
<GID>775</GID>
<name>IN_6</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-42,23.5,-42</points>
<connection>
<GID>697</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>720</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-44.5,24.5,-40</points>
<intersection>-44.5 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-44.5,27.5,-44.5</points>
<connection>
<GID>775</GID>
<name>IN_7</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-40,24.5,-40</points>
<connection>
<GID>696</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>721</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-101.5,27,-98.5</points>
<connection>
<GID>817</GID>
<name>IN_0</name></connection>
<intersection>-101.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-101.5,27,-101.5</points>
<connection>
<GID>725</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>722</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-99.5,26,-97.5</points>
<intersection>-99.5 2</intersection>
<intersection>-97.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-97.5,27,-97.5</points>
<connection>
<GID>817</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-99.5,26,-99.5</points>
<connection>
<GID>713</GID>
<name>IN_0</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>723</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-97.5,24.5,-96.5</points>
<intersection>-97.5 2</intersection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-96.5,27,-96.5</points>
<connection>
<GID>817</GID>
<name>IN_2</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-97.5,24.5,-97.5</points>
<connection>
<GID>710</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>724</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,-95.5,27,-95.5</points>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<connection>
<GID>817</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>725</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-94.5,22,-93.5</points>
<intersection>-94.5 1</intersection>
<intersection>-93.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-94.5,27,-94.5</points>
<connection>
<GID>817</GID>
<name>IN_4</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-93.5,22,-93.5</points>
<connection>
<GID>707</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>726</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-93.5,23.5,-91.5</points>
<intersection>-93.5 1</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-93.5,27,-93.5</points>
<connection>
<GID>817</GID>
<name>IN_5</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-91.5,23.5,-91.5</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>727</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-92.5,24.5,-89.5</points>
<intersection>-92.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-92.5,27,-92.5</points>
<connection>
<GID>817</GID>
<name>IN_6</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-89.5,24.5,-89.5</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>728</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-91.5,25.5,-87.5</points>
<intersection>-91.5 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-91.5,27,-91.5</points>
<connection>
<GID>817</GID>
<name>IN_7</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21.5,-87.5,25.5,-87.5</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>729</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-83.5,147.5,-80</points>
<connection>
<GID>819</GID>
<name>OUT_7</name></connection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>147.5,-80,152,-80</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>730</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-84.5,148.5,-82</points>
<intersection>-84.5 2</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148.5,-82,152,-82</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-84.5,148.5,-84.5</points>
<connection>
<GID>819</GID>
<name>OUT_6</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>731</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-85.5,149.5,-84</points>
<intersection>-85.5 2</intersection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-84,152,-84</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-85.5,149.5,-85.5</points>
<connection>
<GID>819</GID>
<name>OUT_5</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>732</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-86.5,149.5,-86</points>
<intersection>-86.5 2</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-86,152,-86</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-86.5,149.5,-86.5</points>
<connection>
<GID>819</GID>
<name>OUT_4</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>733</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-88,149.5,-87.5</points>
<intersection>-88 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-88,152,-88</points>
<connection>
<GID>766</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-87.5,149.5,-87.5</points>
<connection>
<GID>819</GID>
<name>OUT_3</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>734</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149.5,-90,149.5,-88.5</points>
<intersection>-90 1</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149.5,-90,152,-90</points>
<connection>
<GID>767</GID>
<name>IN_0</name></connection>
<intersection>149.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-88.5,149.5,-88.5</points>
<connection>
<GID>819</GID>
<name>OUT_2</name></connection>
<intersection>149.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>735</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-92,149,-89.5</points>
<intersection>-92 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,-92,152,-92</points>
<connection>
<GID>768</GID>
<name>IN_0</name></connection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-89.5,149,-89.5</points>
<connection>
<GID>819</GID>
<name>OUT_1</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>736</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-94,148,-90.5</points>
<intersection>-94 1</intersection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,-94,152,-94</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-90.5,148,-90.5</points>
<connection>
<GID>819</GID>
<name>OUT_0</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>737</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-79.5,99,-69.5</points>
<intersection>-79.5 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-69.5,99,-69.5</points>
<connection>
<GID>867</GID>
<name>IN_1</name></connection>
<intersection>89.5 3</intersection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97,-79.5,99,-79.5</points>
<connection>
<GID>865</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>89.5,-69.5,89.5,-64.5</points>
<intersection>-69.5 1</intersection>
<intersection>-64.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>89.5,-64.5,91,-64.5</points>
<connection>
<GID>868</GID>
<name>IN_1</name></connection>
<intersection>89.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>738</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-42.5,30.5,-36</points>
<connection>
<GID>775</GID>
<name>load</name></connection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-36,30.5,-36</points>
<connection>
<GID>691</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>739</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-89.5,30,-83.5</points>
<connection>
<GID>817</GID>
<name>load</name></connection>
<intersection>-83.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-83.5,30,-83.5</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>740</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142.5,-81.5,142.5,-78</points>
<connection>
<GID>819</GID>
<name>load</name></connection>
<intersection>-78 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>159,-78,159,-75</points>
<connection>
<GID>693</GID>
<name>IN_0</name></connection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>142.5,-78,159,-78</points>
<intersection>142.5 0</intersection>
<intersection>159 1</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-218.812,79.7914,-113.162,26.3869</PageViewport>
<gate>
<ID>579</ID>
<type>AA_MUX_2x1</type>
<position>-181,48.5</position>
<input>
<ID>IN_0</ID>281 </input>
<input>
<ID>IN_1</ID>280 </input>
<output>
<ID>OUT</ID>899 </output>
<input>
<ID>SEL_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>580</ID>
<type>DA_FROM</type>
<position>-187,47.5</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-3</lparam></gate>
<gate>
<ID>583</ID>
<type>DA_FROM</type>
<position>-187,37.5</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-1</lparam></gate>
<gate>
<ID>393</ID>
<type>DA_FROM</type>
<position>-229,68</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-7</lparam></gate>
<gate>
<ID>592</ID>
<type>DA_FROM</type>
<position>-187,32.5</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-0</lparam></gate>
<gate>
<ID>593</ID>
<type>DA_FROM</type>
<position>-187,42.5</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-2</lparam></gate>
<gate>
<ID>594</ID>
<type>DA_FROM</type>
<position>-187,49.5</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-3</lparam></gate>
<gate>
<ID>595</ID>
<type>DA_FROM</type>
<position>-187,39.5</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-1</lparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>-229,66</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-6</lparam></gate>
<gate>
<ID>596</ID>
<type>DA_FROM</type>
<position>-187,34.5</position>
<input>
<ID>IN_0</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-0</lparam></gate>
<gate>
<ID>403</ID>
<type>DA_FROM</type>
<position>-229,64</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-5</lparam></gate>
<gate>
<ID>597</ID>
<type>DA_FROM</type>
<position>-187,44.5</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-2</lparam></gate>
<gate>
<ID>404</ID>
<type>DA_FROM</type>
<position>-229,62</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-4</lparam></gate>
<gate>
<ID>598</ID>
<type>AA_MUX_2x1</type>
<position>-181,43.5</position>
<input>
<ID>IN_0</ID>283 </input>
<input>
<ID>IN_1</ID>282 </input>
<output>
<ID>OUT</ID>898 </output>
<input>
<ID>SEL_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>405</ID>
<type>DA_FROM</type>
<position>-229,60</position>
<input>
<ID>IN_0</ID>238 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-3</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_SMALL_INVERTER</type>
<position>-223.5,66</position>
<input>
<ID>IN_0</ID>239 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>599</ID>
<type>AA_MUX_2x1</type>
<position>-181,38.5</position>
<input>
<ID>IN_0</ID>286 </input>
<input>
<ID>IN_1</ID>285 </input>
<output>
<ID>OUT</ID>897 </output>
<input>
<ID>SEL_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>DA_FROM</type>
<position>-229,58</position>
<input>
<ID>IN_0</ID>237 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-2</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_MUX_2x1</type>
<position>-181,33.5</position>
<input>
<ID>IN_0</ID>290 </input>
<input>
<ID>IN_1</ID>289 </input>
<output>
<ID>OUT</ID>896 </output>
<input>
<ID>SEL_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>-229,56</position>
<input>
<ID>IN_0</ID>234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-1</lparam></gate>
<gate>
<ID>606</ID>
<type>DE_TO</type>
<position>-158.5,51</position>
<input>
<ID>IN_0</ID>893 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID REG-IS-ZERO</lparam></gate>
<gate>
<ID>413</ID>
<type>DA_FROM</type>
<position>-229,54</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-0</lparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>-224.5,73</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-ADD</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_SMALL_INVERTER</type>
<position>-223.5,64</position>
<input>
<ID>IN_0</ID>241 </input>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>430</ID>
<type>EE_VDD</type>
<position>-214.5,69</position>
<output>
<ID>OUT_0</ID>555 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>627</ID>
<type>BE_NOR4</type>
<position>-175,61</position>
<input>
<ID>IN_0</ID>413 </input>
<input>
<ID>IN_1</ID>412 </input>
<input>
<ID>IN_2</ID>411 </input>
<input>
<ID>IN_3</ID>410 </input>
<output>
<ID>OUT</ID>895 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>50</ID>
<type>AE_REGISTER8</type>
<position>-215.5,60.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>62 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>64 </input>
<input>
<ID>IN_5</ID>65 </input>
<input>
<ID>IN_6</ID>75 </input>
<input>
<ID>IN_7</ID>66 </input>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>41 </output>
<output>
<ID>OUT_2</ID>42 </output>
<output>
<ID>OUT_3</ID>43 </output>
<output>
<ID>OUT_4</ID>44 </output>
<output>
<ID>OUT_5</ID>45 </output>
<output>
<ID>OUT_6</ID>46 </output>
<output>
<ID>OUT_7</ID>40 </output>
<input>
<ID>clock</ID>110 </input>
<input>
<ID>count_enable</ID>242 </input>
<input>
<ID>count_up</ID>555 </input>
<input>
<ID>load</ID>47 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>52</ID>
<type>DE_TO</type>
<position>-207.5,67</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-7</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>-207.5,63</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-5</lparam></gate>
<gate>
<ID>54</ID>
<type>DE_TO</type>
<position>-207.5,61</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-4</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>-207.5,59</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-3</lparam></gate>
<gate>
<ID>56</ID>
<type>DE_TO</type>
<position>-207.5,57</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-2</lparam></gate>
<gate>
<ID>57</ID>
<type>DE_TO</type>
<position>-207.5,55</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-1</lparam></gate>
<gate>
<ID>58</ID>
<type>DE_TO</type>
<position>-207.5,53</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-0</lparam></gate>
<gate>
<ID>59</ID>
<type>DE_TO</type>
<position>-207.5,65</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-6</lparam></gate>
<gate>
<ID>61</ID>
<type>DA_FROM</type>
<position>-224.5,71</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-NEGATOR</lparam></gate>
<gate>
<ID>260</ID>
<type>DA_FROM</type>
<position>-229,50</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CLOCK-PULSE-IN</lparam></gate>
<gate>
<ID>88</ID>
<type>AE_SMALL_INVERTER</type>
<position>-223.5,62</position>
<input>
<ID>IN_0</ID>235 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_SMALL_INVERTER</type>
<position>-223.5,60</position>
<input>
<ID>IN_0</ID>238 </input>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>896</ID>
<type>AA_LABEL</type>
<position>-216,77</position>
<gparam>LABEL_TEXT Negator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1094</ID>
<type>AA_AND2</type>
<position>-165.5,51</position>
<input>
<ID>IN_0</ID>895 </input>
<input>
<ID>IN_1</ID>900 </input>
<output>
<ID>OUT</ID>893 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AE_SMALL_INVERTER</type>
<position>-223.5,58</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1095</ID>
<type>BE_NOR4</type>
<position>-173.5,41.5</position>
<input>
<ID>IN_0</ID>899 </input>
<input>
<ID>IN_1</ID>898 </input>
<input>
<ID>IN_2</ID>897 </input>
<input>
<ID>IN_3</ID>896 </input>
<output>
<ID>OUT</ID>900 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>917</ID>
<type>AA_LABEL</type>
<position>-185,77</position>
<gparam>LABEL_TEXT Comparator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>AE_SMALL_INVERTER</type>
<position>-223.5,56</position>
<input>
<ID>IN_0</ID>234 </input>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>151</ID>
<type>AE_SMALL_INVERTER</type>
<position>-223.5,54</position>
<input>
<ID>IN_0</ID>240 </input>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>152</ID>
<type>AE_SMALL_INVERTER</type>
<position>-223.5,68</position>
<input>
<ID>IN_0</ID>236 </input>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>561</ID>
<type>AA_MUX_2x1</type>
<position>-181,68.5</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>266 </input>
<output>
<ID>OUT</ID>413 </output>
<input>
<ID>SEL_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>562</ID>
<type>DA_FROM</type>
<position>-187,67.5</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-7</lparam></gate>
<gate>
<ID>563</ID>
<type>DA_FROM</type>
<position>-187,57.5</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-5</lparam></gate>
<gate>
<ID>565</ID>
<type>DA_FROM</type>
<position>-187,52.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-4</lparam></gate>
<gate>
<ID>1723</ID>
<type>AA_LABEL</type>
<position>-201.5,80.5</position>
<gparam>LABEL_TEXT Functional Units</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>566</ID>
<type>DA_FROM</type>
<position>-187,62.5</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-6</lparam></gate>
<gate>
<ID>567</ID>
<type>DA_FROM</type>
<position>-187,69.5</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-7</lparam></gate>
<gate>
<ID>568</ID>
<type>DA_FROM</type>
<position>-187,59.5</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-5</lparam></gate>
<gate>
<ID>569</ID>
<type>DA_FROM</type>
<position>-187,54.5</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-4</lparam></gate>
<gate>
<ID>570</ID>
<type>DA_FROM</type>
<position>-187,64.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-6</lparam></gate>
<gate>
<ID>571</ID>
<type>AA_MUX_2x1</type>
<position>-181,63.5</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>269 </input>
<output>
<ID>OUT</ID>412 </output>
<input>
<ID>SEL_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>572</ID>
<type>AA_MUX_2x1</type>
<position>-181,58.5</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>271 </input>
<output>
<ID>OUT</ID>411 </output>
<input>
<ID>SEL_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>573</ID>
<type>AA_MUX_2x1</type>
<position>-181,53.5</position>
<input>
<ID>IN_0</ID>274 </input>
<input>
<ID>IN_1</ID>273 </input>
<output>
<ID>OUT</ID>410 </output>
<input>
<ID>SEL_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>574</ID>
<type>DA_FROM</type>
<position>-187,72.5</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID REG-SELECT</lparam></gate>
<wire>
<ID>410</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-178.5,53.5,-178.5,58</points>
<intersection>53.5 4</intersection>
<intersection>58 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-178.5,58,-178,58</points>
<connection>
<GID>627</GID>
<name>IN_3</name></connection>
<intersection>-178.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-179,53.5,-178.5,53.5</points>
<connection>
<GID>573</GID>
<name>OUT</name></connection>
<intersection>-178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>411</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-178.5,58.5,-178.5,60</points>
<intersection>58.5 3</intersection>
<intersection>60 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-178.5,60,-178,60</points>
<connection>
<GID>627</GID>
<name>IN_2</name></connection>
<intersection>-178.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-179,58.5,-178.5,58.5</points>
<connection>
<GID>572</GID>
<name>OUT</name></connection>
<intersection>-178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>412</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-178.5,62,-178.5,63.5</points>
<intersection>62 2</intersection>
<intersection>63.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-178.5,62,-178,62</points>
<connection>
<GID>627</GID>
<name>IN_1</name></connection>
<intersection>-178.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-179,63.5,-178.5,63.5</points>
<connection>
<GID>571</GID>
<name>OUT</name></connection>
<intersection>-178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-178.5,64,-178.5,68.5</points>
<intersection>64 2</intersection>
<intersection>68.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-178.5,64,-178,64</points>
<connection>
<GID>627</GID>
<name>IN_0</name></connection>
<intersection>-178.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-179,68.5,-178.5,68.5</points>
<connection>
<GID>561</GID>
<name>OUT</name></connection>
<intersection>-178.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-219.5,54,-219.5,57.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>54 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-221.5,54,-219.5,54</points>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection>
<intersection>-219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-211.5,53,-211.5,57.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,53,-209.5,53</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-211.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-211.5,64.5,-211.5,67</points>
<connection>
<GID>50</GID>
<name>OUT_7</name></connection>
<intersection>67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,67,-209.5,67</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-211.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-211,55,-211,58.5</points>
<intersection>55 4</intersection>
<intersection>58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,58.5,-211,58.5</points>
<connection>
<GID>50</GID>
<name>OUT_1</name></connection>
<intersection>-211 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-211,55,-209.5,55</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>-211 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-227,56,-225.5,56</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-210.5,57,-210.5,59.5</points>
<intersection>57 2</intersection>
<intersection>59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,59.5,-210.5,59.5</points>
<connection>
<GID>50</GID>
<name>OUT_2</name></connection>
<intersection>-210.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-210.5,57,-209.5,57</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-210.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-227,62,-225.5,62</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-210,59,-210,60.5</points>
<intersection>59 3</intersection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,60.5,-210,60.5</points>
<connection>
<GID>50</GID>
<name>OUT_3</name></connection>
<intersection>-210 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-210,59,-209.5,59</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-210 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-227,68,-225.5,68</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-210,61,-210,61.5</points>
<intersection>61 3</intersection>
<intersection>61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,61.5,-210,61.5</points>
<connection>
<GID>50</GID>
<name>OUT_4</name></connection>
<intersection>-210 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-210,61,-209.5,61</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-210 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-227,58,-225.5,58</points>
<connection>
<GID>406</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-210,62.5,-210,63</points>
<intersection>62.5 1</intersection>
<intersection>63 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,62.5,-210,62.5</points>
<connection>
<GID>50</GID>
<name>OUT_5</name></connection>
<intersection>-210 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-210,63,-209.5,63</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-210 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-227,60,-225.5,60</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<connection>
<GID>103</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-210,63.5,-210,65</points>
<intersection>63.5 1</intersection>
<intersection>65 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-211.5,63.5,-210,63.5</points>
<connection>
<GID>50</GID>
<name>OUT_6</name></connection>
<intersection>-210 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-210,65,-209.5,65</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-210 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-227,66,-225.5,66</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-216.5,66.5,-216.5,71</points>
<connection>
<GID>50</GID>
<name>load</name></connection>
<intersection>71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-222.5,71,-216.5,71</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-227,54,-225.5,54</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-227,64,-225.5,64</points>
<connection>
<GID>403</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-215.5,66.5,-215.5,73</points>
<connection>
<GID>50</GID>
<name>count_enable</name></connection>
<intersection>73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-222.5,73,-215.5,73</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>-215.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-220,56,-220,58.5</points>
<intersection>56 2</intersection>
<intersection>58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-220,58.5,-219.5,58.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-221.5,56,-220,56</points>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection>
<intersection>-220 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-220.5,58,-220.5,59.5</points>
<intersection>58 3</intersection>
<intersection>59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-220.5,59.5,-219.5,59.5</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>-220.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-221.5,58,-220.5,58</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>-220.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-221,60,-221,60.5</points>
<intersection>60 3</intersection>
<intersection>60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-221,60.5,-219.5,60.5</points>
<connection>
<GID>50</GID>
<name>IN_3</name></connection>
<intersection>-221 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-221.5,60,-221,60</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>-221 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-221,61.5,-221,62</points>
<intersection>61.5 1</intersection>
<intersection>62 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-221,61.5,-219.5,61.5</points>
<connection>
<GID>50</GID>
<name>IN_4</name></connection>
<intersection>-221 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-221.5,62,-221,62</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<intersection>-221 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-220.5,62.5,-220.5,64</points>
<intersection>62.5 1</intersection>
<intersection>64 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-220.5,62.5,-219.5,62.5</points>
<connection>
<GID>50</GID>
<name>IN_5</name></connection>
<intersection>-220.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-221.5,64,-220.5,64</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-220.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-219.5,64.5,-219.5,68</points>
<connection>
<GID>50</GID>
<name>IN_7</name></connection>
<intersection>68 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-221.5,68,-219.5,68</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<intersection>-219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,69.5,-183,69.5</points>
<connection>
<GID>561</GID>
<name>IN_1</name></connection>
<connection>
<GID>567</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,67.5,-183,67.5</points>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<connection>
<GID>562</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-220,63.5,-220,66</points>
<intersection>63.5 1</intersection>
<intersection>66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-220,63.5,-219.5,63.5</points>
<connection>
<GID>50</GID>
<name>IN_6</name></connection>
<intersection>-220 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-221.5,66,-220,66</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>-220 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,64.5,-183,64.5</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<connection>
<GID>571</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,62.5,-183,62.5</points>
<connection>
<GID>566</GID>
<name>IN_0</name></connection>
<connection>
<GID>571</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,59.5,-183,59.5</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<connection>
<GID>572</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,57.5,-183,57.5</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<connection>
<GID>572</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,54.5,-183,54.5</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<connection>
<GID>573</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,52.5,-183,52.5</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<connection>
<GID>573</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-184,36,-184,72.5</points>
<intersection>36 25</intersection>
<intersection>41 28</intersection>
<intersection>46 27</intersection>
<intersection>51 26</intersection>
<intersection>56 5</intersection>
<intersection>61 6</intersection>
<intersection>66 7</intersection>
<intersection>71 1</intersection>
<intersection>72.5 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-184,71,-181,71</points>
<connection>
<GID>561</GID>
<name>SEL_0</name></connection>
<intersection>-184 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-184,56,-181,56</points>
<connection>
<GID>573</GID>
<name>SEL_0</name></connection>
<intersection>-184 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-184,61,-181,61</points>
<connection>
<GID>572</GID>
<name>SEL_0</name></connection>
<intersection>-184 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-184,66,-181,66</points>
<connection>
<GID>571</GID>
<name>SEL_0</name></connection>
<intersection>-184 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-185,72.5,-184,72.5</points>
<connection>
<GID>574</GID>
<name>IN_0</name></connection>
<intersection>-184 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-184,36,-181,36</points>
<connection>
<GID>600</GID>
<name>SEL_0</name></connection>
<intersection>-184 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-184,51,-181,51</points>
<connection>
<GID>579</GID>
<name>SEL_0</name></connection>
<intersection>-184 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-184,46,-181,46</points>
<connection>
<GID>598</GID>
<name>SEL_0</name></connection>
<intersection>-184 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-184,41,-181,41</points>
<connection>
<GID>599</GID>
<name>SEL_0</name></connection>
<intersection>-184 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,49.5,-183,49.5</points>
<connection>
<GID>579</GID>
<name>IN_1</name></connection>
<connection>
<GID>594</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,47.5,-183,47.5</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<connection>
<GID>580</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,44.5,-183,44.5</points>
<connection>
<GID>597</GID>
<name>IN_0</name></connection>
<connection>
<GID>598</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,42.5,-183,42.5</points>
<connection>
<GID>593</GID>
<name>IN_0</name></connection>
<connection>
<GID>598</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,39.5,-183,39.5</points>
<connection>
<GID>595</GID>
<name>IN_0</name></connection>
<connection>
<GID>599</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,37.5,-183,37.5</points>
<connection>
<GID>583</GID>
<name>IN_0</name></connection>
<connection>
<GID>599</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,34.5,-183,34.5</points>
<connection>
<GID>596</GID>
<name>IN_0</name></connection>
<connection>
<GID>600</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-185,32.5,-183,32.5</points>
<connection>
<GID>592</GID>
<name>IN_0</name></connection>
<connection>
<GID>600</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-216.5,50,-216.5,55.5</points>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-227,50,-216.5,50</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>-216.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>893</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-162.5,51,-160.5,51</points>
<connection>
<GID>606</GID>
<name>IN_0</name></connection>
<connection>
<GID>1094</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>895</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-169.5,52,-169.5,61</points>
<intersection>52 2</intersection>
<intersection>61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-171,61,-169.5,61</points>
<connection>
<GID>627</GID>
<name>OUT</name></connection>
<intersection>-169.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-169.5,52,-168.5,52</points>
<connection>
<GID>1094</GID>
<name>IN_0</name></connection>
<intersection>-169.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>896</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-176.5,33.5,-176.5,38.5</points>
<connection>
<GID>1095</GID>
<name>IN_3</name></connection>
<intersection>33.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-179,33.5,-176.5,33.5</points>
<connection>
<GID>600</GID>
<name>OUT</name></connection>
<intersection>-176.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>897</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-177.5,38.5,-177.5,40.5</points>
<intersection>38.5 1</intersection>
<intersection>40.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-179,38.5,-177.5,38.5</points>
<connection>
<GID>599</GID>
<name>OUT</name></connection>
<intersection>-177.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-177.5,40.5,-176.5,40.5</points>
<connection>
<GID>1095</GID>
<name>IN_2</name></connection>
<intersection>-177.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>898</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-177.5,42.5,-177.5,43.5</points>
<intersection>42.5 2</intersection>
<intersection>43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-179,43.5,-177.5,43.5</points>
<connection>
<GID>598</GID>
<name>OUT</name></connection>
<intersection>-177.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-177.5,42.5,-176.5,42.5</points>
<connection>
<GID>1095</GID>
<name>IN_1</name></connection>
<intersection>-177.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>899</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-177.5,44.5,-177.5,48.5</points>
<intersection>44.5 2</intersection>
<intersection>48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-179,48.5,-177.5,48.5</points>
<connection>
<GID>579</GID>
<name>OUT</name></connection>
<intersection>-177.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-177.5,44.5,-176.5,44.5</points>
<connection>
<GID>1095</GID>
<name>IN_0</name></connection>
<intersection>-177.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>900</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-169,41.5,-169,50</points>
<intersection>41.5 2</intersection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-169,50,-168.5,50</points>
<connection>
<GID>1094</GID>
<name>IN_1</name></connection>
<intersection>-169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-169.5,41.5,-169,41.5</points>
<connection>
<GID>1095</GID>
<name>OUT</name></connection>
<intersection>-169 0</intersection></hsegment></shape></wire>
<wire>
<ID>555</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-214.5,66.5,-214.5,68</points>
<connection>
<GID>50</GID>
<name>count_up</name></connection>
<connection>
<GID>430</GID>
<name>OUT_0</name></connection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>-212.365,154.095,13.3679,39.99</PageViewport>
<gate>
<ID>193</ID>
<type>DE_TO</type>
<position>-148,69.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-0</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_MUX_2x1</type>
<position>-153,84.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>104 </output>
<input>
<ID>SEL_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>195</ID>
<type>DA_FROM</type>
<position>-159,83.5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-3</lparam></gate>
<gate>
<ID>196</ID>
<type>DA_FROM</type>
<position>-159,73.5</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-1</lparam></gate>
<gate>
<ID>197</ID>
<type>DA_FROM</type>
<position>-159,68.5</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-0</lparam></gate>
<gate>
<ID>391</ID>
<type>DA_FROM</type>
<position>-75.5,110</position>
<input>
<ID>IN_0</ID>599 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID USE-USER-INSTRUCTION</lparam></gate>
<gate>
<ID>198</ID>
<type>DA_FROM</type>
<position>-159,78.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-2</lparam></gate>
<gate>
<ID>199</ID>
<type>DA_FROM</type>
<position>-159,85.5</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-3</lparam></gate>
<gate>
<ID>200</ID>
<type>DA_FROM</type>
<position>-159,75.5</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-1</lparam></gate>
<gate>
<ID>779</ID>
<type>AA_MUX_2x1</type>
<position>-78,77</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>830 </output>
<input>
<ID>SEL_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>DA_FROM</type>
<position>-159,70.5</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-0</lparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>-159,80.5</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-2</lparam></gate>
<gate>
<ID>781</ID>
<type>DE_TO</type>
<position>-59.5,83.5</position>
<input>
<ID>IN_0</ID>834 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-RAM-1</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_MUX_2x1</type>
<position>-153,79.5</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>105 </output>
<input>
<ID>SEL_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_MUX_2x1</type>
<position>-153,74.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>106 </output>
<input>
<ID>SEL_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_MUX_2x1</type>
<position>-153,69.5</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>107 </output>
<input>
<ID>SEL_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_MUX_2x1</type>
<position>-194.5,73.5</position>
<input>
<ID>IN_0</ID>170 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>175 </output>
<input>
<ID>SEL_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>DA_FROM</type>
<position>-206,75.5</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-3</lparam></gate>
<gate>
<ID>787</ID>
<type>DA_FROM</type>
<position>-84,87.5</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-USER-2</lparam></gate>
<gate>
<ID>209</ID>
<type>DE_TO</type>
<position>-189,96.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-IN-6</lparam></gate>
<gate>
<ID>210</ID>
<type>DE_TO</type>
<position>-189,88.5</position>
<input>
<ID>IN_0</ID>164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-IN-5</lparam></gate>
<gate>
<ID>983</ID>
<type>DA_FROM</type>
<position>-71,100.5</position>
<input>
<ID>IN_0</ID>823 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID RUN-PROGRAM</lparam></gate>
<gate>
<ID>211</ID>
<type>DE_TO</type>
<position>-189.5,81</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-IN-4</lparam></gate>
<gate>
<ID>212</ID>
<type>DE_TO</type>
<position>-189.5,73.5</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-IN-3</lparam></gate>
<gate>
<ID>791</ID>
<type>DA_FROM</type>
<position>-84,93.5</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-USER-3</lparam></gate>
<gate>
<ID>213</ID>
<type>DE_TO</type>
<position>-189.5,65.5</position>
<input>
<ID>IN_0</ID>224 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-IN-2</lparam></gate>
<gate>
<ID>792</ID>
<type>DA_FROM</type>
<position>-84,76</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-USER-0</lparam></gate>
<gate>
<ID>214</ID>
<type>DE_TO</type>
<position>-189.5,58</position>
<input>
<ID>IN_0</ID>250 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-IN-1</lparam></gate>
<gate>
<ID>215</ID>
<type>DE_TO</type>
<position>-189,50</position>
<input>
<ID>IN_0</ID>353 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-IN-0</lparam></gate>
<gate>
<ID>794</ID>
<type>DA_FROM</type>
<position>-84,81.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-USER-1</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_MUX_2x1</type>
<position>-200.5,72.5</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>174 </input>
<output>
<ID>OUT</ID>170 </output>
<input>
<ID>SEL_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>795</ID>
<type>DE_TO</type>
<position>-59.5,78</position>
<input>
<ID>IN_0</ID>835 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-RAM-0</lparam></gate>
<gate>
<ID>989</ID>
<type>DA_FROM</type>
<position>-70,90.5</position>
<input>
<ID>IN_0</ID>828 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-2</lparam></gate>
<gate>
<ID>217</ID>
<type>DA_FROM</type>
<position>-206,71.5</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-3</lparam></gate>
<gate>
<ID>990</ID>
<type>DA_FROM</type>
<position>-70,79</position>
<input>
<ID>IN_0</ID>831 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-0</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>-206,65.5</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-2</lparam></gate>
<gate>
<ID>797</ID>
<type>AA_LABEL</type>
<position>-72.5,114</position>
<gparam>LABEL_TEXT IR RAM Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>991</ID>
<type>DA_FROM</type>
<position>-70,96.5</position>
<input>
<ID>IN_0</ID>825 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-3</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_MUX_2x1</type>
<position>-194.5,65.5</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>177 </input>
<output>
<ID>OUT</ID>224 </output>
<input>
<ID>SEL_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>992</ID>
<type>DA_FROM</type>
<position>-70,84.5</position>
<input>
<ID>IN_0</ID>829 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-1</lparam></gate>
<gate>
<ID>220</ID>
<type>DA_FROM</type>
<position>-206,67.5</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-2</lparam></gate>
<gate>
<ID>993</ID>
<type>AA_MUX_2x1</type>
<position>-66,89.5</position>
<input>
<ID>IN_0</ID>826 </input>
<input>
<ID>IN_1</ID>828 </input>
<output>
<ID>OUT</ID>833 </output>
<input>
<ID>SEL_0</ID>823 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_MUX_2x1</type>
<position>-200.5,64.5</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>179 </input>
<output>
<ID>OUT</ID>176 </output>
<input>
<ID>SEL_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>994</ID>
<type>AA_MUX_2x1</type>
<position>-66,83.5</position>
<input>
<ID>IN_0</ID>827 </input>
<input>
<ID>IN_1</ID>829 </input>
<output>
<ID>OUT</ID>834 </output>
<input>
<ID>SEL_0</ID>823 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>-206,63.5</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-2</lparam></gate>
<gate>
<ID>995</ID>
<type>AA_MUX_2x1</type>
<position>-66,78</position>
<input>
<ID>IN_0</ID>830 </input>
<input>
<ID>IN_1</ID>831 </input>
<output>
<ID>OUT</ID>835 </output>
<input>
<ID>SEL_0</ID>823 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>223</ID>
<type>DA_FROM</type>
<position>-206,58</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-1</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_MUX_2x1</type>
<position>-194.5,58</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>247 </input>
<output>
<ID>OUT</ID>250 </output>
<input>
<ID>SEL_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>997</ID>
<type>AA_LABEL</type>
<position>-157.5,114.5</position>
<gparam>LABEL_TEXT R0 Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>DA_FROM</type>
<position>-206,60</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-1</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_MUX_2x1</type>
<position>-200.5,57</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>245 </output>
<input>
<ID>SEL_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>-206,56</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-1</lparam></gate>
<gate>
<ID>236</ID>
<type>DA_FROM</type>
<position>-205.5,50</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-0</lparam></gate>
<gate>
<ID>237</ID>
<type>AA_MUX_2x1</type>
<position>-194,50</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>353 </output>
<input>
<ID>SEL_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>431</ID>
<type>DE_TO</type>
<position>-60,104</position>
<input>
<ID>IN_0</ID>600 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READY-TO-SAVE-INSTRUCTION</lparam></gate>
<gate>
<ID>238</ID>
<type>DA_FROM</type>
<position>-205.5,52</position>
<input>
<ID>IN_0</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-0</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_MUX_2x1</type>
<position>-200,49</position>
<input>
<ID>IN_0</ID>253 </input>
<input>
<ID>IN_1</ID>254 </input>
<output>
<ID>OUT</ID>251 </output>
<input>
<ID>SEL_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>DA_FROM</type>
<position>-205.5,48</position>
<input>
<ID>IN_0</ID>253 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-0</lparam></gate>
<gate>
<ID>436</ID>
<type>DA_FROM</type>
<position>-121,86</position>
<input>
<ID>IN_0</ID>501 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-3</lparam></gate>
<gate>
<ID>437</ID>
<type>DA_FROM</type>
<position>-121,76</position>
<input>
<ID>IN_0</ID>502 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-1</lparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>-121,71</position>
<input>
<ID>IN_0</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-0</lparam></gate>
<gate>
<ID>448</ID>
<type>DA_FROM</type>
<position>-121,81</position>
<input>
<ID>IN_0</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-2</lparam></gate>
<gate>
<ID>449</ID>
<type>DA_FROM</type>
<position>-121,106</position>
<input>
<ID>IN_0</ID>519 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-7</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>-205.5,104</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-7</lparam></gate>
<gate>
<ID>450</ID>
<type>DA_FROM</type>
<position>-121,96</position>
<input>
<ID>IN_0</ID>529 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-5</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>-121,91</position>
<input>
<ID>IN_0</ID>526 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-4</lparam></gate>
<gate>
<ID>452</ID>
<type>DA_FROM</type>
<position>-121,101</position>
<input>
<ID>IN_0</ID>527 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-6</lparam></gate>
<gate>
<ID>1043</ID>
<type>AA_LABEL</type>
<position>-117.5,114.5</position>
<gparam>LABEL_TEXT R1 Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>853</ID>
<type>AA_MUX_2x1</type>
<position>-66,95.5</position>
<input>
<ID>IN_0</ID>824 </input>
<input>
<ID>IN_1</ID>825 </input>
<output>
<ID>OUT</ID>832 </output>
<input>
<ID>SEL_0</ID>823 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>673</ID>
<type>AE_OR2</type>
<position>-159,109.5</position>
<input>
<ID>IN_0</ID>605 </input>
<input>
<ID>IN_1</ID>604 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_MUX_2x1</type>
<position>-194,104</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>131 </input>
<output>
<ID>OUT</ID>133 </output>
<input>
<ID>SEL_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>DA_FROM</type>
<position>-214.5,108</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID REG-SELECT</lparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>-205.5,106</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-7</lparam></gate>
<gate>
<ID>509</ID>
<type>AA_AND2</type>
<position>-66.5,104</position>
<input>
<ID>IN_0</ID>597 </input>
<input>
<ID>IN_1</ID>602 </input>
<output>
<ID>OUT</ID>600 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>DE_TO</type>
<position>-189,104</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-IN-7</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>-214.5,111</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID LOAD-IN</lparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>-205.5,96.5</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-6</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_MUX_2x1</type>
<position>-194,96.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>155 </output>
<input>
<ID>SEL_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>709</ID>
<type>DA_FROM</type>
<position>-128,111</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID OP-SUB</lparam></gate>
<gate>
<ID>1096</ID>
<type>AA_LABEL</type>
<position>-199,114.5</position>
<gparam>LABEL_TEXT MBR Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>DA_FROM</type>
<position>-205.5,98.5</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-6</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_MUX_2x1</type>
<position>-200,95.5</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>134 </output>
<input>
<ID>SEL_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>DA_FROM</type>
<position>-205.5,94.5</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-6</lparam></gate>
<gate>
<ID>714</ID>
<type>DA_FROM</type>
<position>-165.5,110.5</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID OP-SUB</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>-205.5,88.5</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-5</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_MUX_2x1</type>
<position>-194,88.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>164 </output>
<input>
<ID>SEL_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>-205.5,90.5</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-5</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_MUX_2x1</type>
<position>-200,87.5</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>156 </output>
<input>
<ID>SEL_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>-205.5,86.5</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-5</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>-206,81</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-4</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_MUX_2x1</type>
<position>-194.5,81</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>169 </output>
<input>
<ID>SEL_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>721</ID>
<type>AE_OR2</type>
<position>-121.5,110</position>
<input>
<ID>IN_0</ID>607 </input>
<input>
<ID>IN_1</ID>606 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>-206,83</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IN-4</lparam></gate>
<gate>
<ID>337</ID>
<type>DA_FROM</type>
<position>-75.5,108</position>
<input>
<ID>IN_0</ID>597 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID WRITE-INSTRUCTION</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_MUX_2x1</type>
<position>-200.5,80</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>168 </input>
<output>
<ID>OUT</ID>165 </output>
<input>
<ID>SEL_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>730</ID>
<type>AE_SMALL_INVERTER</type>
<position>-73,103</position>
<input>
<ID>IN_0</ID>528 </input>
<output>
<ID>OUT_0</ID>602 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>345</ID>
<type>DE_TO</type>
<position>-110,70</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-0</lparam></gate>
<gate>
<ID>346</ID>
<type>AA_MUX_2x1</type>
<position>-115,85</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>501 </input>
<output>
<ID>OUT</ID>221 </output>
<input>
<ID>SEL_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>DA_FROM</type>
<position>-206,79</position>
<input>
<ID>IN_0</ID>167 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-4</lparam></gate>
<gate>
<ID>732</ID>
<type>DA_FROM</type>
<position>-84,89.5</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-2</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>-121,84</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-3</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>-206,73.5</position>
<input>
<ID>IN_0</ID>174 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-3</lparam></gate>
<gate>
<ID>733</ID>
<type>DA_FROM</type>
<position>-84,95.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-3</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_MUX_2x1</type>
<position>-200,103</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>130 </output>
<input>
<ID>SEL_0</ID>161 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>-121,74</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-1</lparam></gate>
<gate>
<ID>734</ID>
<type>DA_FROM</type>
<position>-84,78</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-0</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>-205.5,102</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-7</lparam></gate>
<gate>
<ID>349</ID>
<type>DA_FROM</type>
<position>-121,69</position>
<input>
<ID>IN_0</ID>217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-0</lparam></gate>
<gate>
<ID>735</ID>
<type>DA_FROM</type>
<position>-84,83.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MAR-1</lparam></gate>
<gate>
<ID>350</ID>
<type>DA_FROM</type>
<position>-121,79</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-2</lparam></gate>
<gate>
<ID>737</ID>
<type>AA_MUX_2x1</type>
<position>-78,94.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>824 </output>
<input>
<ID>SEL_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>738</ID>
<type>AA_MUX_2x1</type>
<position>-78,88.5</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>826 </output>
<input>
<ID>SEL_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>739</ID>
<type>DE_TO</type>
<position>-59.5,89.5</position>
<input>
<ID>IN_0</ID>833 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-RAM-2</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_MUX_2x1</type>
<position>-115,80</position>
<input>
<ID>IN_0</ID>205 </input>
<input>
<ID>IN_1</ID>503 </input>
<output>
<ID>OUT</ID>222 </output>
<input>
<ID>SEL_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_MUX_2x1</type>
<position>-115,75</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>223 </output>
<input>
<ID>SEL_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_MUX_2x1</type>
<position>-115,70</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>506 </input>
<output>
<ID>OUT</ID>246 </output>
<input>
<ID>SEL_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_MUX_2x1</type>
<position>-115,105</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>519 </input>
<output>
<ID>OUT</ID>220 </output>
<input>
<ID>SEL_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>-121,104</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-7</lparam></gate>
<gate>
<ID>360</ID>
<type>DA_FROM</type>
<position>-121,94</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-5</lparam></gate>
<gate>
<ID>361</ID>
<type>DA_FROM</type>
<position>-121,89</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-4</lparam></gate>
<gate>
<ID>362</ID>
<type>DA_FROM</type>
<position>-121,99</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-6</lparam></gate>
<gate>
<ID>748</ID>
<type>DE_TO</type>
<position>-59.5,95.5</position>
<input>
<ID>IN_0</ID>832 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-RAM-3</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_MUX_2x1</type>
<position>-153,104.5</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>103 </output>
<input>
<ID>SEL_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_SMALL_INVERTER</type>
<position>-82.5,108</position>
<input>
<ID>IN_0</ID>597 </input>
<output>
<ID>OUT_0</ID>598 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>-159,103.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-7</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_MUX_2x1</type>
<position>-115,100</position>
<input>
<ID>IN_0</ID>196 </input>
<input>
<ID>IN_1</ID>527 </input>
<output>
<ID>OUT</ID>218 </output>
<input>
<ID>SEL_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>-159,93.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-5</lparam></gate>
<gate>
<ID>368</ID>
<type>AA_MUX_2x1</type>
<position>-115,95</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>529 </input>
<output>
<ID>OUT</ID>219 </output>
<input>
<ID>SEL_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>-159,88.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-4</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_MUX_2x1</type>
<position>-115,90</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>526 </input>
<output>
<ID>OUT</ID>225 </output>
<input>
<ID>SEL_0</ID>201 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>-159,98.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-6</lparam></gate>
<gate>
<ID>1720</ID>
<type>AA_LABEL</type>
<position>-158,119.5</position>
<gparam>LABEL_TEXT Busses</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>-159,105.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-7</lparam></gate>
<gate>
<ID>756</ID>
<type>AA_MUX_2x1</type>
<position>-78,82.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>71 </input>
<output>
<ID>OUT</ID>827 </output>
<input>
<ID>SEL_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>DA_FROM</type>
<position>-159,95.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-5</lparam></gate>
<gate>
<ID>372</ID>
<type>DA_FROM</type>
<position>-128,109</position>
<input>
<ID>IN_0</ID>606 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID OP-ADD</lparam></gate>
<gate>
<ID>179</ID>
<type>DA_FROM</type>
<position>-159,90.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-4</lparam></gate>
<gate>
<ID>373</ID>
<type>DE_TO</type>
<position>-110,105</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-7</lparam></gate>
<gate>
<ID>180</ID>
<type>DA_FROM</type>
<position>-159,100.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-6</lparam></gate>
<gate>
<ID>374</ID>
<type>DE_TO</type>
<position>-110,100</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-6</lparam></gate>
<gate>
<ID>181</ID>
<type>AA_MUX_2x1</type>
<position>-153,99.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>101 </output>
<input>
<ID>SEL_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>DE_TO</type>
<position>-110,95</position>
<input>
<ID>IN_0</ID>219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-5</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_MUX_2x1</type>
<position>-153,94.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>102 </output>
<input>
<ID>SEL_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>DE_TO</type>
<position>-110,90</position>
<input>
<ID>IN_0</ID>225 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-4</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_MUX_2x1</type>
<position>-153,89.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>108 </output>
<input>
<ID>SEL_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>DE_TO</type>
<position>-110,85</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-3</lparam></gate>
<gate>
<ID>378</ID>
<type>DE_TO</type>
<position>-110,80</position>
<input>
<ID>IN_0</ID>222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-2</lparam></gate>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>-165.5,108.5</position>
<input>
<ID>IN_0</ID>604 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID OP-ADD</lparam></gate>
<gate>
<ID>379</ID>
<type>DE_TO</type>
<position>-110,75</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-IN-1</lparam></gate>
<gate>
<ID>186</ID>
<type>DE_TO</type>
<position>-148,104.5</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-7</lparam></gate>
<gate>
<ID>187</ID>
<type>DE_TO</type>
<position>-148,99.5</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-6</lparam></gate>
<gate>
<ID>188</ID>
<type>DE_TO</type>
<position>-148,94.5</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-5</lparam></gate>
<gate>
<ID>189</ID>
<type>DE_TO</type>
<position>-148,89.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-4</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_TO</type>
<position>-148,84.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-3</lparam></gate>
<gate>
<ID>384</ID>
<type>AA_AND2</type>
<position>-82.5,103</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>599 </input>
<output>
<ID>OUT</ID>528 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>DE_TO</type>
<position>-148,79.5</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-2</lparam></gate>
<gate>
<ID>192</ID>
<type>DE_TO</type>
<position>-148,74.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-IN-1</lparam></gate>
<wire>
<ID>194</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,104,-117,104</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<connection>
<GID>359</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,99,-117,99</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,94,-117,94</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,89,-117,89</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<connection>
<GID>369</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-118,72.5,-118,110</points>
<intersection>72.5 20</intersection>
<intersection>77.5 21</intersection>
<intersection>82.5 22</intersection>
<intersection>87.5 23</intersection>
<intersection>92.5 5</intersection>
<intersection>97.5 6</intersection>
<intersection>102.5 7</intersection>
<intersection>107.5 1</intersection>
<intersection>110 40</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-118,107.5,-115,107.5</points>
<connection>
<GID>358</GID>
<name>SEL_0</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-118,92.5,-115,92.5</points>
<connection>
<GID>369</GID>
<name>SEL_0</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-118,97.5,-115,97.5</points>
<connection>
<GID>368</GID>
<name>SEL_0</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-118,102.5,-115,102.5</points>
<connection>
<GID>367</GID>
<name>SEL_0</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-118,72.5,-115,72.5</points>
<connection>
<GID>357</GID>
<name>SEL_0</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-118,77.5,-115,77.5</points>
<connection>
<GID>356</GID>
<name>SEL_0</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-118,82.5,-115,82.5</points>
<connection>
<GID>355</GID>
<name>SEL_0</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-118,87.5,-115,87.5</points>
<connection>
<GID>346</GID>
<name>SEL_0</name></connection>
<intersection>-118 0</intersection></hsegment>
<hsegment>
<ID>40</ID>
<points>-118.5,110,-118,110</points>
<connection>
<GID>721</GID>
<name>OUT</name></connection>
<intersection>-118 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,84,-117,84</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<connection>
<GID>347</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,79,-117,79</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<connection>
<GID>355</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,74,-117,74</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>356</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>597</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-80.5,105,-80.5,108</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>105 1</intersection>
<intersection>108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-80.5,105,-69.5,105</points>
<connection>
<GID>509</GID>
<name>IN_0</name></connection>
<intersection>-80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-80.5,108,-77.5,108</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>-80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>598</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-86.5,104,-86.5,108</points>
<intersection>104 3</intersection>
<intersection>108 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-86.5,108,-84.5,108</points>
<connection>
<GID>366</GID>
<name>OUT_0</name></connection>
<intersection>-86.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-86.5,104,-85.5,104</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>-86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>599</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,102,-87.5,110</points>
<intersection>102 1</intersection>
<intersection>110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-87.5,102,-85.5,102</points>
<connection>
<GID>384</GID>
<name>IN_1</name></connection>
<intersection>-87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-87.5,110,-77.5,110</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>-87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>600</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-63.5,104,-62,104</points>
<connection>
<GID>509</GID>
<name>OUT</name></connection>
<connection>
<GID>431</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>602</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-71,103,-69.5,103</points>
<connection>
<GID>730</GID>
<name>OUT_0</name></connection>
<connection>
<GID>509</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,69,-117,69</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<connection>
<GID>357</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,100,-112,100</points>
<connection>
<GID>367</GID>
<name>OUT</name></connection>
<connection>
<GID>374</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>604</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-163.5,108.5,-162,108.5</points>
<connection>
<GID>673</GID>
<name>IN_1</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,95,-112,95</points>
<connection>
<GID>368</GID>
<name>OUT</name></connection>
<connection>
<GID>375</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>605</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-163.5,110.5,-162,110.5</points>
<connection>
<GID>673</GID>
<name>IN_0</name></connection>
<connection>
<GID>714</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,105,-112,105</points>
<connection>
<GID>358</GID>
<name>OUT</name></connection>
<connection>
<GID>373</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>606</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-126,109,-124.5,109</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<connection>
<GID>721</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,85,-112,85</points>
<connection>
<GID>346</GID>
<name>OUT</name></connection>
<connection>
<GID>377</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>607</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-126,111,-124.5,111</points>
<connection>
<GID>721</GID>
<name>IN_0</name></connection>
<connection>
<GID>709</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,80,-112,80</points>
<connection>
<GID>355</GID>
<name>OUT</name></connection>
<connection>
<GID>378</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,75,-112,75</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<connection>
<GID>379</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-192.5,65.5,-191.5,65.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<connection>
<GID>219</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,90,-112,90</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<connection>
<GID>376</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>823</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74,98,-74,100.5</points>
<intersection>98 2</intersection>
<intersection>100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74,100.5,-73,100.5</points>
<connection>
<GID>983</GID>
<name>IN_0</name></connection>
<intersection>-74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-74,98,-62.5,98</points>
<connection>
<GID>853</GID>
<name>SEL_0</name></connection>
<intersection>-74 0</intersection>
<intersection>-62.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-62.5,80.5,-62.5,98</points>
<intersection>80.5 8</intersection>
<intersection>86 9</intersection>
<intersection>92 10</intersection>
<intersection>98 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-66,80.5,-62.5,80.5</points>
<connection>
<GID>995</GID>
<name>SEL_0</name></connection>
<intersection>-62.5 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-66,86,-62.5,86</points>
<connection>
<GID>994</GID>
<name>SEL_0</name></connection>
<intersection>-62.5 4</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-66,92,-62.5,92</points>
<connection>
<GID>993</GID>
<name>SEL_0</name></connection>
<intersection>-62.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>824</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76,94.5,-68,94.5</points>
<connection>
<GID>737</GID>
<name>OUT</name></connection>
<connection>
<GID>853</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-198.5,57,-196.5,57</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>226</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>825</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-68,96.5,-68,96.5</points>
<connection>
<GID>853</GID>
<name>IN_1</name></connection>
<connection>
<GID>991</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113,70,-112,70</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>357</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>826</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76,88.5,-68,88.5</points>
<connection>
<GID>738</GID>
<name>OUT</name></connection>
<connection>
<GID>993</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,60,-199.5,60</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-199.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-199.5,59,-199.5,60</points>
<intersection>59 9</intersection>
<intersection>60 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-199.5,59,-196.5,59</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>-199.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>827</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76,82.5,-68,82.5</points>
<connection>
<GID>756</GID>
<name>OUT</name></connection>
<connection>
<GID>994</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,76,-80,76</points>
<connection>
<GID>792</GID>
<name>IN_0</name></connection>
<connection>
<GID>779</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,56,-202.5,56</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<connection>
<GID>227</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>828</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-68,90.5,-68,90.5</points>
<connection>
<GID>989</GID>
<name>IN_0</name></connection>
<connection>
<GID>993</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,58,-202.5,58</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<connection>
<GID>226</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>829</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-68,84.5,-68,84.5</points>
<connection>
<GID>992</GID>
<name>IN_0</name></connection>
<connection>
<GID>994</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,78,-80,78</points>
<connection>
<GID>734</GID>
<name>IN_0</name></connection>
<connection>
<GID>779</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-192.5,58,-191.5,58</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<connection>
<GID>224</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>830</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76,77,-68,77</points>
<connection>
<GID>779</GID>
<name>OUT</name></connection>
<connection>
<GID>995</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-198,49,-196,49</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<connection>
<GID>239</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>831</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68,79,-68,79</points>
<connection>
<GID>990</GID>
<name>IN_0</name></connection>
<connection>
<GID>995</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,52,-199,52</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>-199 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-199,51,-199,52</points>
<intersection>51 9</intersection>
<intersection>52 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-199,51,-196,51</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<intersection>-199 8</intersection></hsegment></shape></wire>
<wire>
<ID>832</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,95.5,-61.5,95.5</points>
<connection>
<GID>853</GID>
<name>OUT</name></connection>
<connection>
<GID>748</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,48,-202,48</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<connection>
<GID>240</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>833</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,89.5,-61.5,89.5</points>
<connection>
<GID>993</GID>
<name>OUT</name></connection>
<connection>
<GID>739</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-203.5,50,-202,50</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<connection>
<GID>239</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>834</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,83.5,-61.5,83.5</points>
<connection>
<GID>994</GID>
<name>OUT</name></connection>
<connection>
<GID>781</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>835</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,78,-61.5,78</points>
<connection>
<GID>995</GID>
<name>OUT</name></connection>
<connection>
<GID>795</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,93.5,-80,93.5</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<connection>
<GID>791</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,81.5,-80,81.5</points>
<connection>
<GID>756</GID>
<name>IN_0</name></connection>
<connection>
<GID>794</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,87.5,-80,87.5</points>
<connection>
<GID>738</GID>
<name>IN_0</name></connection>
<connection>
<GID>787</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,83.5,-80,83.5</points>
<connection>
<GID>756</GID>
<name>IN_1</name></connection>
<connection>
<GID>735</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,95.5,-80,95.5</points>
<connection>
<GID>737</GID>
<name>IN_1</name></connection>
<connection>
<GID>733</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-82,89.5,-80,89.5</points>
<connection>
<GID>738</GID>
<name>IN_1</name></connection>
<connection>
<GID>732</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,105.5,-155,105.5</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<connection>
<GID>177</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,103.5,-155,103.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<connection>
<GID>173</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,100.5,-155,100.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<connection>
<GID>181</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,98.5,-155,98.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<connection>
<GID>181</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,95.5,-155,95.5</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<connection>
<GID>182</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,93.5,-155,93.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<connection>
<GID>182</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,90.5,-155,90.5</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<connection>
<GID>183</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,88.5,-155,88.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<connection>
<GID>183</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-156,72,-156,109.5</points>
<connection>
<GID>673</GID>
<name>OUT</name></connection>
<intersection>72 20</intersection>
<intersection>77 21</intersection>
<intersection>82 22</intersection>
<intersection>87 23</intersection>
<intersection>92 5</intersection>
<intersection>97 6</intersection>
<intersection>102 7</intersection>
<intersection>107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-156,107,-153,107</points>
<connection>
<GID>172</GID>
<name>SEL_0</name></connection>
<intersection>-156 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-156,92,-153,92</points>
<connection>
<GID>183</GID>
<name>SEL_0</name></connection>
<intersection>-156 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-156,97,-153,97</points>
<connection>
<GID>182</GID>
<name>SEL_0</name></connection>
<intersection>-156 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-156,102,-153,102</points>
<connection>
<GID>181</GID>
<name>SEL_0</name></connection>
<intersection>-156 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-156,72,-153,72</points>
<connection>
<GID>205</GID>
<name>SEL_0</name></connection>
<intersection>-156 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-156,77,-153,77</points>
<connection>
<GID>204</GID>
<name>SEL_0</name></connection>
<intersection>-156 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-156,82,-153,82</points>
<connection>
<GID>203</GID>
<name>SEL_0</name></connection>
<intersection>-156 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-156,87,-153,87</points>
<connection>
<GID>194</GID>
<name>SEL_0</name></connection>
<intersection>-156 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,85.5,-155,85.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<connection>
<GID>199</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,83.5,-155,83.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<connection>
<GID>195</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,80.5,-155,80.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<connection>
<GID>203</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,78.5,-155,78.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<connection>
<GID>203</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,75.5,-155,75.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<connection>
<GID>204</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,73.5,-155,73.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<connection>
<GID>204</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,70.5,-155,70.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>205</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-157,68.5,-155,68.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<connection>
<GID>205</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-151,99.5,-150,99.5</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<connection>
<GID>187</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-151,94.5,-150,94.5</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<connection>
<GID>188</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-151,104.5,-150,104.5</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-151,84.5,-150,84.5</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<connection>
<GID>190</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-151,79.5,-150,79.5</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<connection>
<GID>191</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-151,74.5,-150,74.5</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<connection>
<GID>192</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-151,69.5,-150,69.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<connection>
<GID>205</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-151,89.5,-150,89.5</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>501</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,86,-117,86</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>346</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>502</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,76,-117,76</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<connection>
<GID>356</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>503</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,81,-117,81</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<connection>
<GID>355</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>506</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,71,-117,71</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<connection>
<GID>357</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-198,103,-196,103</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,106,-199,106</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-199 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-199,105,-199,106</points>
<intersection>105 9</intersection>
<intersection>106 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-199,105,-196,105</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>-199 8</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-192,104,-191,104</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>519</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,106,-117,106</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<connection>
<GID>358</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-198,95.5,-196,95.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,98.5,-199,98.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-199 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-199,97.5,-199,98.5</points>
<intersection>97.5 9</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-199,97.5,-196,97.5</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>-199 8</intersection></hsegment></shape></wire>
<wire>
<ID>526</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,91,-117,91</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<connection>
<GID>369</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>527</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,101,-117,101</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,94.5,-202,94.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>528</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81,79.5,-81,97</points>
<intersection>79.5 4</intersection>
<intersection>85 3</intersection>
<intersection>91 5</intersection>
<intersection>97 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-81,97,-78,97</points>
<intersection>-81 0</intersection>
<intersection>-78 36</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-81,85,-78,85</points>
<connection>
<GID>756</GID>
<name>SEL_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-81,79.5,-78,79.5</points>
<connection>
<GID>779</GID>
<name>SEL_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-81,91,-78,91</points>
<connection>
<GID>738</GID>
<name>SEL_0</name></connection>
<intersection>-81 0</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>-78,97,-78,103</points>
<connection>
<GID>737</GID>
<name>SEL_0</name></connection>
<intersection>97 2</intersection>
<intersection>103 37</intersection></vsegment>
<hsegment>
<ID>37</ID>
<points>-79.5,103,-75,103</points>
<connection>
<GID>384</GID>
<name>OUT</name></connection>
<connection>
<GID>730</GID>
<name>IN_0</name></connection>
<intersection>-78 36</intersection></hsegment></shape></wire>
<wire>
<ID>529</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,96,-117,96</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,96.5,-202,96.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-197,54,-197,111</points>
<intersection>54 19</intersection>
<intersection>62 20</intersection>
<intersection>69.5 21</intersection>
<intersection>77.5 22</intersection>
<intersection>84.5 23</intersection>
<intersection>92.5 13</intersection>
<intersection>100 3</intersection>
<intersection>108 4</intersection>
<intersection>111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212.5,111,-197,111</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-197 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-197,100,-194,100</points>
<intersection>-197 0</intersection>
<intersection>-194 8</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-197,108,-194,108</points>
<intersection>-197 0</intersection>
<intersection>-194 29</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-194,99,-194,100</points>
<connection>
<GID>128</GID>
<name>SEL_0</name></connection>
<intersection>100 3</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-197,92.5,-194,92.5</points>
<intersection>-197 0</intersection>
<intersection>-194 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-194,91,-194,92.5</points>
<connection>
<GID>136</GID>
<name>SEL_0</name></connection>
<intersection>92.5 13</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-197,54,-194,54</points>
<intersection>-197 0</intersection>
<intersection>-194 28</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-197,62,-194.5,62</points>
<intersection>-197 0</intersection>
<intersection>-194.5 27</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-197,69.5,-194.5,69.5</points>
<intersection>-197 0</intersection>
<intersection>-194.5 26</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-197,77.5,-194.5,77.5</points>
<intersection>-197 0</intersection>
<intersection>-194.5 25</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-197,84.5,-194.5,84.5</points>
<intersection>-197 0</intersection>
<intersection>-194.5 24</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>-194.5,83.5,-194.5,84.5</points>
<connection>
<GID>141</GID>
<name>SEL_0</name></connection>
<intersection>84.5 23</intersection></vsegment>
<vsegment>
<ID>25</ID>
<points>-194.5,76,-194.5,77.5</points>
<connection>
<GID>207</GID>
<name>SEL_0</name></connection>
<intersection>77.5 22</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>-194.5,68,-194.5,69.5</points>
<connection>
<GID>219</GID>
<name>SEL_0</name></connection>
<intersection>69.5 21</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>-194.5,60.5,-194.5,62</points>
<connection>
<GID>224</GID>
<name>SEL_0</name></connection>
<intersection>62 20</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>-194,52.5,-194,54</points>
<connection>
<GID>237</GID>
<name>SEL_0</name></connection>
<intersection>54 19</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>-194,106.5,-194,108</points>
<connection>
<GID>116</GID>
<name>SEL_0</name></connection>
<intersection>108 4</intersection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-192,96.5,-191,96.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<connection>
<GID>128</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-198,87.5,-196,87.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,102,-202,102</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>156</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,104,-202,104</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,90.5,-199,90.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-199 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-199,89.5,-199,90.5</points>
<intersection>89.5 9</intersection>
<intersection>90.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-199,89.5,-196,89.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>-199 8</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,86.5,-202,86.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>353</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-192,50,-191,50</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<connection>
<GID>237</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-212.5,53.5,-212.5,108</points>
<intersection>53.5 24</intersection>
<intersection>61.5 25</intersection>
<intersection>69 26</intersection>
<intersection>77 27</intersection>
<intersection>84.5 28</intersection>
<intersection>92 18</intersection>
<intersection>100 12</intersection>
<intersection>108 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-212.5,108,-200,108</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-212.5 0</intersection>
<intersection>-200 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-200,105.5,-200,108</points>
<connection>
<GID>155</GID>
<name>SEL_0</name></connection>
<intersection>108 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-212.5,100,-200,100</points>
<intersection>-212.5 0</intersection>
<intersection>-200 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-200,98,-200,100</points>
<connection>
<GID>133</GID>
<name>SEL_0</name></connection>
<intersection>100 12</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-212.5,92,-200,92</points>
<intersection>-212.5 0</intersection>
<intersection>-200 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-200,90,-200,92</points>
<connection>
<GID>138</GID>
<name>SEL_0</name></connection>
<intersection>92 18</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-212.5,53.5,-200,53.5</points>
<intersection>-212.5 0</intersection>
<intersection>-200 33</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>-212.5,61.5,-200.5,61.5</points>
<intersection>-212.5 0</intersection>
<intersection>-200.5 32</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-212.5,69,-200.5,69</points>
<intersection>-212.5 0</intersection>
<intersection>-200.5 31</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-212.5,77,-200.5,77</points>
<intersection>-212.5 0</intersection>
<intersection>-200.5 30</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-212.5,84.5,-200.5,84.5</points>
<intersection>-212.5 0</intersection>
<intersection>-200.5 29</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>-200.5,82.5,-200.5,84.5</points>
<connection>
<GID>148</GID>
<name>SEL_0</name></connection>
<intersection>84.5 28</intersection></vsegment>
<vsegment>
<ID>30</ID>
<points>-200.5,75,-200.5,77</points>
<connection>
<GID>216</GID>
<name>SEL_0</name></connection>
<intersection>77 27</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>-200.5,67,-200.5,69</points>
<connection>
<GID>221</GID>
<name>SEL_0</name></connection>
<intersection>69 26</intersection></vsegment>
<vsegment>
<ID>32</ID>
<points>-200.5,59.5,-200.5,61.5</points>
<connection>
<GID>226</GID>
<name>SEL_0</name></connection>
<intersection>61.5 25</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>-200,51.5,-200,53.5</points>
<connection>
<GID>239</GID>
<name>SEL_0</name></connection>
<intersection>53.5 24</intersection></vsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-203.5,88.5,-202,88.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-192,88.5,-191,88.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-198.5,80,-196.5,80</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,83,-199.5,83</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-199.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-199.5,82,-199.5,83</points>
<intersection>82 9</intersection>
<intersection>83 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-199.5,82,-196.5,82</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>-199.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,79,-202.5,79</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<connection>
<GID>153</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,81,-202.5,81</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-192.5,81,-191.5,81</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>141</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-198.5,72.5,-196.5,72.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>216</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,75.5,-199.5,75.5</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>-199.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-199.5,74.5,-199.5,75.5</points>
<intersection>74.5 9</intersection>
<intersection>75.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-199.5,74.5,-196.5,74.5</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<intersection>-199.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,71.5,-202.5,71.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<connection>
<GID>217</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,73.5,-202.5,73.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<connection>
<GID>154</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-192.5,73.5,-191.5,73.5</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<connection>
<GID>212</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-198.5,64.5,-196.5,64.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<connection>
<GID>221</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,67.5,-199.5,67.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>-199.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-199.5,66.5,-199.5,67.5</points>
<intersection>66.5 9</intersection>
<intersection>67.5 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-199.5,66.5,-196.5,66.5</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>-199.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,63.5,-202.5,63.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<connection>
<GID>222</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-204,65.5,-202.5,65.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>221</GID>
<name>IN_1</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-212.896,6.09055,-73.0537,-64.5981</PageViewport>
<gate>
<ID>206</ID>
<type>DA_FROM</type>
<position>-174.5,-34.5</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-4</lparam></gate>
<gate>
<ID>1561</ID>
<type>AA_LABEL</type>
<position>-167,-8</position>
<gparam>LABEL_TEXT Adder Op 1 Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1597</ID>
<type>AA_LABEL</type>
<position>-120,-7.5</position>
<gparam>LABEL_TEXT Adder Op 2 Bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>-174.5,-24.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-6</lparam></gate>
<gate>
<ID>248</ID>
<type>DA_FROM</type>
<position>-174.5,-17.5</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-7</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>-174.5,-27.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-5</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>-174.5,-32.5</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-4</lparam></gate>
<gate>
<ID>251</ID>
<type>DA_FROM</type>
<position>-174.5,-22.5</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-6</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_MUX_2x1</type>
<position>-168.5,-23.5</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>346 </output>
<input>
<ID>SEL_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_MUX_2x1</type>
<position>-168.5,-28.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>347 </output>
<input>
<ID>SEL_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_MUX_2x1</type>
<position>-168.5,-33.5</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>348 </output>
<input>
<ID>SEL_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>DA_FROM</type>
<position>-174.5,-14.5</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID OP-SUB</lparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>-126.5,-33.5</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-4</lparam></gate>
<gate>
<ID>268</ID>
<type>DA_FROM</type>
<position>-126.5,-23.5</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-6</lparam></gate>
<gate>
<ID>269</ID>
<type>DA_FROM</type>
<position>-126.5,-16.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-7</lparam></gate>
<gate>
<ID>270</ID>
<type>DA_FROM</type>
<position>-126.5,-26.5</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-5</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>-126.5,-31.5</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-4</lparam></gate>
<gate>
<ID>272</ID>
<type>DA_FROM</type>
<position>-126.5,-21.5</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-6</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_MUX_2x1</type>
<position>-120.5,-22.5</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>258 </input>
<output>
<ID>OUT</ID>297 </output>
<input>
<ID>SEL_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>AA_MUX_2x1</type>
<position>-120.5,-27.5</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>260 </input>
<output>
<ID>OUT</ID>298 </output>
<input>
<ID>SEL_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>275</ID>
<type>AA_MUX_2x1</type>
<position>-120.5,-32.5</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>262 </input>
<output>
<ID>OUT</ID>328 </output>
<input>
<ID>SEL_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>292</ID>
<type>DA_FROM</type>
<position>-126.5,-13.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID REG-SELECT</lparam></gate>
<gate>
<ID>293</ID>
<type>DE_TO</type>
<position>-115.5,-17.5</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-7</lparam></gate>
<gate>
<ID>294</ID>
<type>DE_TO</type>
<position>-115.5,-22.5</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-6</lparam></gate>
<gate>
<ID>295</ID>
<type>DE_TO</type>
<position>-115.5,-27.5</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-5</lparam></gate>
<gate>
<ID>296</ID>
<type>DE_TO</type>
<position>-115.5,-32.5</position>
<input>
<ID>IN_0</ID>328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-4</lparam></gate>
<gate>
<ID>297</ID>
<type>DE_TO</type>
<position>-115.5,-37.5</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-3</lparam></gate>
<gate>
<ID>298</ID>
<type>DE_TO</type>
<position>-115.5,-42.5</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-2</lparam></gate>
<gate>
<ID>299</ID>
<type>DE_TO</type>
<position>-115.5,-47.5</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-1</lparam></gate>
<gate>
<ID>300</ID>
<type>DE_TO</type>
<position>-115.5,-52.5</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-2-0</lparam></gate>
<gate>
<ID>301</ID>
<type>AA_MUX_2x1</type>
<position>-120.5,-37.5</position>
<input>
<ID>IN_0</ID>276 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>300 </output>
<input>
<ID>SEL_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>DA_FROM</type>
<position>-126.5,-38.5</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-3</lparam></gate>
<gate>
<ID>303</ID>
<type>DA_FROM</type>
<position>-126.5,-48.5</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-1</lparam></gate>
<gate>
<ID>304</ID>
<type>DA_FROM</type>
<position>-126.5,-53.5</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-0</lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>-126.5,-43.5</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-2</lparam></gate>
<gate>
<ID>306</ID>
<type>DA_FROM</type>
<position>-126.5,-36.5</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-3</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>-126.5,-46.5</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-1</lparam></gate>
<gate>
<ID>308</ID>
<type>DA_FROM</type>
<position>-126.5,-51.5</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-0</lparam></gate>
<gate>
<ID>309</ID>
<type>DA_FROM</type>
<position>-126.5,-41.5</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R1-2</lparam></gate>
<gate>
<ID>310</ID>
<type>AA_MUX_2x1</type>
<position>-120.5,-42.5</position>
<input>
<ID>IN_0</ID>278 </input>
<input>
<ID>IN_1</ID>277 </input>
<output>
<ID>OUT</ID>301 </output>
<input>
<ID>SEL_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>AA_MUX_2x1</type>
<position>-120.5,-47.5</position>
<input>
<ID>IN_0</ID>331 </input>
<input>
<ID>IN_1</ID>279 </input>
<output>
<ID>OUT</ID>302 </output>
<input>
<ID>SEL_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>312</ID>
<type>AA_MUX_2x1</type>
<position>-120.5,-52.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>295 </input>
<output>
<ID>OUT</ID>303 </output>
<input>
<ID>SEL_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>313</ID>
<type>AA_MUX_2x1</type>
<position>-120.5,-17.5</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>256 </input>
<output>
<ID>OUT</ID>299 </output>
<input>
<ID>SEL_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>-126.5,-18.5</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-7</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>-126.5,-28.5</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R0-5</lparam></gate>
<gate>
<ID>316</ID>
<type>DE_TO</type>
<position>-163.5,-18.5</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-7</lparam></gate>
<gate>
<ID>317</ID>
<type>DE_TO</type>
<position>-163.5,-23.5</position>
<input>
<ID>IN_0</ID>346 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-6</lparam></gate>
<gate>
<ID>318</ID>
<type>DE_TO</type>
<position>-163.5,-28.5</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-5</lparam></gate>
<gate>
<ID>319</ID>
<type>DE_TO</type>
<position>-163.5,-33.5</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-4</lparam></gate>
<gate>
<ID>320</ID>
<type>DE_TO</type>
<position>-163.5,-38.5</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-3</lparam></gate>
<gate>
<ID>321</ID>
<type>DE_TO</type>
<position>-163.5,-43.5</position>
<input>
<ID>IN_0</ID>351 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-2</lparam></gate>
<gate>
<ID>322</ID>
<type>DE_TO</type>
<position>-163.5,-48.5</position>
<input>
<ID>IN_0</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-1</lparam></gate>
<gate>
<ID>323</ID>
<type>DE_TO</type>
<position>-163.5,-53.5</position>
<input>
<ID>IN_0</ID>345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-IN-1-0</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_MUX_2x1</type>
<position>-168.5,-38.5</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>188 </input>
<output>
<ID>OUT</ID>350 </output>
<input>
<ID>SEL_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>-174.5,-39.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-3</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>-174.5,-49.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-1</lparam></gate>
<gate>
<ID>160</ID>
<type>DA_FROM</type>
<position>-174.5,-54.5</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-0</lparam></gate>
<gate>
<ID>161</ID>
<type>DA_FROM</type>
<position>-174.5,-44.5</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-2</lparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>-174.5,-37.5</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-3</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>-174.5,-47.5</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-1</lparam></gate>
<gate>
<ID>164</ID>
<type>DA_FROM</type>
<position>-174.5,-52.5</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-0</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>-174.5,-42.5</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-2</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_MUX_2x1</type>
<position>-168.5,-43.5</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>351 </output>
<input>
<ID>SEL_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_MUX_2x1</type>
<position>-168.5,-48.5</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>344 </output>
<input>
<ID>SEL_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_MUX_2x1</type>
<position>-168.5,-53.5</position>
<input>
<ID>IN_0</ID>244 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>345 </output>
<input>
<ID>SEL_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_MUX_2x1</type>
<position>-168.5,-18.5</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>349 </output>
<input>
<ID>SEL_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>DA_FROM</type>
<position>-174.5,-19.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-7</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>-174.5,-29.5</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MBR-5</lparam></gate>
<gate>
<ID>1721</ID>
<type>AA_LABEL</type>
<position>-141,-3.5</position>
<gparam>LABEL_TEXT Busses</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-52.5,-170.5,-52.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-54.5,-170.5,-54.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-49.5,-170.5,-49.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<connection>
<GID>159</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-16.5,-122.5,-16.5</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124.5,-18.5,-122.5,-18.5</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<connection>
<GID>314</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-21.5,-122.5,-21.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<connection>
<GID>272</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-23.5,-122.5,-23.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<connection>
<GID>268</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-26.5,-122.5,-26.5</points>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<connection>
<GID>270</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124.5,-28.5,-122.5,-28.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<connection>
<GID>315</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-31.5,-122.5,-31.5</points>
<connection>
<GID>275</GID>
<name>IN_1</name></connection>
<connection>
<GID>271</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-33.5,-122.5,-33.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<connection>
<GID>267</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-123.5,-50,-123.5,-13.5</points>
<intersection>-50 20</intersection>
<intersection>-45 21</intersection>
<intersection>-40 22</intersection>
<intersection>-35 23</intersection>
<intersection>-30 5</intersection>
<intersection>-25 6</intersection>
<intersection>-20 7</intersection>
<intersection>-15 1</intersection>
<intersection>-13.5 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-123.5,-15,-120.5,-15</points>
<connection>
<GID>313</GID>
<name>SEL_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-123.5,-30,-120.5,-30</points>
<connection>
<GID>275</GID>
<name>SEL_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-123.5,-25,-120.5,-25</points>
<connection>
<GID>274</GID>
<name>SEL_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-123.5,-20,-120.5,-20</points>
<connection>
<GID>273</GID>
<name>SEL_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-124.5,-13.5,-123.5,-13.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-123.5,-50,-120.5,-50</points>
<connection>
<GID>312</GID>
<name>SEL_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-123.5,-45,-120.5,-45</points>
<connection>
<GID>311</GID>
<name>SEL_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-123.5,-40,-120.5,-40</points>
<connection>
<GID>310</GID>
<name>SEL_0</name></connection>
<intersection>-123.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-123.5,-35,-120.5,-35</points>
<connection>
<GID>301</GID>
<name>SEL_0</name></connection>
<intersection>-123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124.5,-36.5,-122.5,-36.5</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<connection>
<GID>306</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124.5,-38.5,-122.5,-38.5</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-41.5,-122.5,-41.5</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<connection>
<GID>309</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-43.5,-122.5,-43.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<connection>
<GID>305</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-46.5,-122.5,-46.5</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<connection>
<GID>307</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-51.5,-122.5,-51.5</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<connection>
<GID>308</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-53.5,-122.5,-53.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<connection>
<GID>304</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-22.5,-117.5,-22.5</points>
<connection>
<GID>273</GID>
<name>OUT</name></connection>
<connection>
<GID>294</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-27.5,-117.5,-27.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<connection>
<GID>295</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-17.5,-117.5,-17.5</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<connection>
<GID>293</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-37.5,-117.5,-37.5</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<connection>
<GID>297</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-42.5,-117.5,-42.5</points>
<connection>
<GID>310</GID>
<name>OUT</name></connection>
<connection>
<GID>298</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-47.5,-117.5,-47.5</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<connection>
<GID>299</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-52.5,-117.5,-52.5</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<connection>
<GID>300</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-118.5,-32.5,-117.5,-32.5</points>
<connection>
<GID>275</GID>
<name>OUT</name></connection>
<connection>
<GID>296</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>331</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-124.5,-48.5,-122.5,-48.5</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<connection>
<GID>303</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>344</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-48.5,-165.5,-48.5</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<connection>
<GID>322</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>345</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-53.5,-165.5,-53.5</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<connection>
<GID>323</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>346</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-23.5,-165.5,-23.5</points>
<connection>
<GID>252</GID>
<name>OUT</name></connection>
<connection>
<GID>317</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>347</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-28.5,-165.5,-28.5</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<connection>
<GID>318</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>348</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-33.5,-165.5,-33.5</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<connection>
<GID>319</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>349</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-18.5,-165.5,-18.5</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<connection>
<GID>316</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>350</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-38.5,-165.5,-38.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<connection>
<GID>320</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>351</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-166.5,-43.5,-165.5,-43.5</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<connection>
<GID>321</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-17.5,-170.5,-17.5</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<connection>
<GID>248</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-19.5,-170.5,-19.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<connection>
<GID>169</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-22.5,-170.5,-22.5</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<connection>
<GID>251</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-24.5,-170.5,-24.5</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<connection>
<GID>247</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-27.5,-170.5,-27.5</points>
<connection>
<GID>253</GID>
<name>IN_1</name></connection>
<connection>
<GID>249</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-29.5,-170.5,-29.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<connection>
<GID>253</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-32.5,-170.5,-32.5</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-34.5,-170.5,-34.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<connection>
<GID>206</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-171.5,-51,-171.5,-14.5</points>
<intersection>-51 20</intersection>
<intersection>-46 21</intersection>
<intersection>-41 22</intersection>
<intersection>-36 23</intersection>
<intersection>-31 5</intersection>
<intersection>-26 6</intersection>
<intersection>-21 7</intersection>
<intersection>-16 1</intersection>
<intersection>-14.5 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-171.5,-16,-168.5,-16</points>
<connection>
<GID>169</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-171.5,-31,-168.5,-31</points>
<connection>
<GID>254</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-171.5,-26,-168.5,-26</points>
<connection>
<GID>253</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-171.5,-21,-168.5,-21</points>
<connection>
<GID>252</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-172.5,-14.5,-171.5,-14.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>-171.5 0</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>-171.5,-51,-168.5,-51</points>
<connection>
<GID>168</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-171.5,-46,-168.5,-46</points>
<connection>
<GID>167</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-171.5,-41,-168.5,-41</points>
<connection>
<GID>166</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-171.5,-36,-168.5,-36</points>
<connection>
<GID>157</GID>
<name>SEL_0</name></connection>
<intersection>-171.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-37.5,-170.5,-37.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<connection>
<GID>162</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-39.5,-170.5,-39.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-42.5,-170.5,-42.5</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<connection>
<GID>165</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-44.5,-170.5,-44.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-172.5,-47.5,-170.5,-47.5</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<connection>
<GID>163</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>-257.435,142.874,-130.265,78.5915</PageViewport>
<gate>
<ID>1</ID>
<type>DA_FROM</type>
<position>-205.5,106</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-DECODE</lparam></gate>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>-179.5,109.5</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-MAR</lparam></gate>
<gate>
<ID>3</ID>
<type>DE_TO</type>
<position>-201.5,103.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-OP</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>-201.5,101</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-REG</lparam></gate>
<gate>
<ID>7</ID>
<type>DA_FROM</type>
<position>-205.5,109.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-FETCH-2</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>-201.5,109.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-IR</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>-205.5,113</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-FETCH-1</lparam></gate>
<gate>
<ID>1316</ID>
<type>AA_LABEL</type>
<position>-198.5,121</position>
<gparam>LABEL_TEXT Command Sequencing</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>380</ID>
<type>AE_OR2</type>
<position>-186,109.5</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-203.5,101,-203.5,106</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-203.5,106,-190.5,106</points>
<intersection>-203.5 0</intersection>
<intersection>-190.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-190.5,106,-190.5,108.5</points>
<intersection>106 1</intersection>
<intersection>108.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-190.5,108.5,-189,108.5</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>-190.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-203.5,109.5,-203.5,109.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-183,109.5,-181.5,109.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>380</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-190.5,110.5,-190.5,113</points>
<intersection>110.5 2</intersection>
<intersection>113 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-203.5,113,-190.5,113</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-190.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-190.5,110.5,-189,110.5</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>-190.5 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>-204.843,117.956,31.0927,-1.30606</PageViewport>
<gate>
<ID>774</ID>
<type>AA_AND2</type>
<position>-85,-45.5</position>
<input>
<ID>IN_0</ID>637 </input>
<input>
<ID>IN_1</ID>585 </input>
<output>
<ID>OUT</ID>584 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>778</ID>
<type>DA_FROM</type>
<position>-78.5,-41.5</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID REG-IS-ZERO</lparam></gate>
<gate>
<ID>782</ID>
<type>DE_TO</type>
<position>-78.5,-45.5</position>
<input>
<ID>IN_0</ID>584 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-PC</lparam></gate>
<gate>
<ID>601</ID>
<type>DA_FROM</type>
<position>-66,14</position>
<input>
<ID>IN_0</ID>464 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-SUB</lparam></gate>
<gate>
<ID>602</ID>
<type>DE_TO</type>
<position>-54.5,75</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OUTPUT-READY</lparam></gate>
<gate>
<ID>604</ID>
<type>DA_FROM</type>
<position>-125.5,89.5</position>
<input>
<ID>IN_0</ID>477 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-READ</lparam></gate>
<gate>
<ID>605</ID>
<type>DA_FROM</type>
<position>-126,80.5</position>
<input>
<ID>IN_0</ID>479 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-2</lparam></gate>
<gate>
<ID>608</ID>
<type>DA_FROM</type>
<position>-125.5,75.5</position>
<input>
<ID>IN_0</ID>480 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-3</lparam></gate>
<gate>
<ID>803</ID>
<type>AE_SMALL_INVERTER</type>
<position>-85,-41.5</position>
<input>
<ID>IN_0</ID>636 </input>
<output>
<ID>OUT_0</ID>637 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>611</ID>
<type>DA_FROM</type>
<position>-125.5,85.5</position>
<input>
<ID>IN_0</ID>478 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-1</lparam></gate>
<gate>
<ID>612</ID>
<type>AA_AND2</type>
<position>-118,86.5</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>478 </input>
<output>
<ID>OUT</ID>483 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>613</ID>
<type>AA_AND2</type>
<position>-61,80.5</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>490 </input>
<output>
<ID>OUT</ID>451 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>614</ID>
<type>AA_AND2</type>
<position>-61,75</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>491 </input>
<output>
<ID>OUT</ID>452 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>615</ID>
<type>AA_AND2</type>
<position>-118,81.5</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>479 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>616</ID>
<type>AA_AND2</type>
<position>-118,76.5</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>480 </input>
<output>
<ID>OUT</ID>379 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>618</ID>
<type>DA_FROM</type>
<position>-131,49.5</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-LOAD</lparam></gate>
<gate>
<ID>619</ID>
<type>DA_FROM</type>
<position>-131.5,40.5</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-2</lparam></gate>
<gate>
<ID>626</ID>
<type>DA_FROM</type>
<position>-131,45.5</position>
<input>
<ID>IN_0</ID>496 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-1</lparam></gate>
<gate>
<ID>242</ID>
<type>DE_TO</type>
<position>-54.5,85.5</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WRITE-LOAD-MBR</lparam></gate>
<gate>
<ID>628</ID>
<type>AA_AND2</type>
<position>-123.5,46.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>496 </input>
<output>
<ID>OUT</ID>453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND2</type>
<position>-61,70</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>429 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>DE_TO</type>
<position>-104,-15</position>
<input>
<ID>IN_0</ID>460 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-R0</lparam></gate>
<gate>
<ID>631</ID>
<type>AA_AND2</type>
<position>-123.5,41.5</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>497 </input>
<output>
<ID>OUT</ID>518 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>DE_TO</type>
<position>-104,-10.5</position>
<input>
<ID>IN_0</ID>457 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-R1</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>-114,-6.5</position>
<input>
<ID>IN_0</ID>458 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID REG-SELECT</lparam></gate>
<gate>
<ID>637</ID>
<type>DA_FROM</type>
<position>-66.5,5</position>
<input>
<ID>IN_0</ID>466 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-2</lparam></gate>
<gate>
<ID>639</ID>
<type>DE_TO</type>
<position>-52,11</position>
<input>
<ID>IN_0</ID>504 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-MBR</lparam></gate>
<gate>
<ID>640</ID>
<type>DA_FROM</type>
<position>-66.5,-0.5</position>
<input>
<ID>IN_0</ID>467 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-3</lparam></gate>
<gate>
<ID>641</ID>
<type>DA_FROM</type>
<position>-66.5,-5.5</position>
<input>
<ID>IN_0</ID>468 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-4</lparam></gate>
<gate>
<ID>642</ID>
<type>DA_FROM</type>
<position>-66.5,-10.5</position>
<input>
<ID>IN_0</ID>469 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-5</lparam></gate>
<gate>
<ID>643</ID>
<type>DA_FROM</type>
<position>-67,-24.5</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-6</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_AND2</type>
<position>-110.5,-10.5</position>
<input>
<ID>IN_0</ID>458 </input>
<input>
<ID>IN_1</ID>459 </input>
<output>
<ID>OUT</ID>457 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>644</ID>
<type>DA_FROM</type>
<position>-67,-29</position>
<input>
<ID>IN_0</ID>471 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-7</lparam></gate>
<gate>
<ID>258</ID>
<type>AE_SMALL_INVERTER</type>
<position>-116.5,-10.5</position>
<input>
<ID>IN_0</ID>458 </input>
<output>
<ID>OUT_0</ID>461 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1031</ID>
<type>DE_TO</type>
<position>-102,90</position>
<input>
<ID>IN_0</ID>857 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STOP-EXECUTION</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_TO</type>
<position>-116.5,46.5</position>
<input>
<ID>IN_0</ID>453 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-LOAD-MBR</lparam></gate>
<gate>
<ID>645</ID>
<type>DA_FROM</type>
<position>-66,10</position>
<input>
<ID>IN_0</ID>465 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-1</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_AND2</type>
<position>-110.5,-15</position>
<input>
<ID>IN_0</ID>461 </input>
<input>
<ID>IN_1</ID>459 </input>
<output>
<ID>OUT</ID>460 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>646</ID>
<type>AA_AND2</type>
<position>-58.5,11</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>465 </input>
<output>
<ID>OUT</ID>504 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1033</ID>
<type>AA_AND2</type>
<position>-109,90</position>
<input>
<ID>IN_0</ID>858 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>857 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>261</ID>
<type>DE_TO</type>
<position>-54,70</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WRITE-SEQ-RESET</lparam></gate>
<gate>
<ID>647</ID>
<type>AA_AND2</type>
<position>-58.5,6</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>466 </input>
<output>
<ID>OUT</ID>505 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>648</ID>
<type>AA_AND2</type>
<position>-58.5,0.5</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>556 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1035</ID>
<type>DA_FROM</type>
<position>-107.5,93.5</position>
<input>
<ID>IN_0</ID>858 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID RUN-PROGRAM</lparam></gate>
<gate>
<ID>263</ID>
<type>DA_FROM</type>
<position>-69,69</position>
<input>
<ID>IN_0</ID>416 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-4</lparam></gate>
<gate>
<ID>649</ID>
<type>AA_AND2</type>
<position>-58.5,-4.5</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>468 </input>
<output>
<ID>OUT</ID>540 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>650</ID>
<type>AA_AND2</type>
<position>-58.5,-9.5</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>469 </input>
<output>
<ID>OUT</ID>537 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>-119.5,97.5</position>
<gparam>LABEL_TEXT Read</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>651</ID>
<type>AA_AND2</type>
<position>-59,-23.5</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>470 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>-62,97.5</position>
<gparam>LABEL_TEXT Write</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>459</ID>
<type>DA_FROM</type>
<position>-126,63.5</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-5</lparam></gate>
<gate>
<ID>652</ID>
<type>AA_AND2</type>
<position>-59,-28</position>
<input>
<ID>IN_0</ID>464 </input>
<input>
<ID>IN_1</ID>471 </input>
<output>
<ID>OUT</ID>608 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>AA_LABEL</type>
<position>-120.5,53.5</position>
<gparam>LABEL_TEXT Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>653</ID>
<type>DA_FROM</type>
<position>-130.5,12</position>
<input>
<ID>IN_0</ID>472 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-ADD</lparam></gate>
<gate>
<ID>654</ID>
<type>DA_FROM</type>
<position>-131,3</position>
<input>
<ID>IN_0</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-2</lparam></gate>
<gate>
<ID>655</ID>
<type>DA_FROM</type>
<position>-131,-2.5</position>
<input>
<ID>IN_0</ID>475 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-3</lparam></gate>
<gate>
<ID>463</ID>
<type>AA_AND2</type>
<position>-118,64.5</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>564 </input>
<output>
<ID>OUT</ID>565 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>656</ID>
<type>DA_FROM</type>
<position>-130.5,8</position>
<input>
<ID>IN_0</ID>473 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-1</lparam></gate>
<gate>
<ID>657</ID>
<type>AA_AND2</type>
<position>-123,9</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>473 </input>
<output>
<ID>OUT</ID>500 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>658</ID>
<type>AA_AND2</type>
<position>-123,4</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>-131.5,28</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-3</lparam></gate>
<gate>
<ID>659</ID>
<type>AA_AND2</type>
<position>-123,-1.5</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>475 </input>
<output>
<ID>OUT</ID>415 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>660</ID>
<type>DE_TO</type>
<position>-116,-1.5</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-ADDER-RESULT</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>-123.5,29</position>
<input>
<ID>IN_0</ID>495 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>661</ID>
<type>DE_TO</type>
<position>-106.5,33</position>
<input>
<ID>IN_0</ID>520 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-LOAD-R0</lparam></gate>
<gate>
<ID>83</ID>
<type>DE_TO</type>
<position>-117,29</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-SEQ-RESET</lparam></gate>
<gate>
<ID>662</ID>
<type>DE_TO</type>
<position>-106.5,37.5</position>
<input>
<ID>IN_0</ID>516 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-LOAD-R1</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>-126,70.5</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-4</lparam></gate>
<gate>
<ID>663</ID>
<type>DE_TO</type>
<position>-116,4</position>
<input>
<ID>IN_0</ID>414 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-ADDER</lparam></gate>
<gate>
<ID>664</ID>
<type>DE_TO</type>
<position>-52,6</position>
<input>
<ID>IN_0</ID>505 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-NEGATOR</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND2</type>
<position>-118,71.5</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>576 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>665</ID>
<type>DE_TO</type>
<position>-51.5,0.5</position>
<input>
<ID>IN_0</ID>556 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NEG-ADD</lparam></gate>
<gate>
<ID>666</ID>
<type>DA_FROM</type>
<position>-116.5,41.5</position>
<input>
<ID>IN_0</ID>517 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID REG-SELECT</lparam></gate>
<gate>
<ID>668</ID>
<type>AA_AND2</type>
<position>-123,-7</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>494 </input>
<output>
<ID>OUT</ID>459 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>-131,-8</position>
<input>
<ID>IN_0</ID>494 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-4</lparam></gate>
<gate>
<ID>670</ID>
<type>AA_AND2</type>
<position>-123,-20</position>
<input>
<ID>IN_0</ID>472 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>462 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>671</ID>
<type>DA_FROM</type>
<position>-131,-21</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-5</lparam></gate>
<gate>
<ID>672</ID>
<type>AA_AND2</type>
<position>-113,37.5</position>
<input>
<ID>IN_0</ID>517 </input>
<input>
<ID>IN_1</ID>518 </input>
<output>
<ID>OUT</ID>516 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>674</ID>
<type>AE_SMALL_INVERTER</type>
<position>-119,37.5</position>
<input>
<ID>IN_0</ID>517 </input>
<output>
<ID>OUT_0</ID>521 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>675</ID>
<type>AA_AND2</type>
<position>-113,33</position>
<input>
<ID>IN_0</ID>521 </input>
<input>
<ID>IN_1</ID>518 </input>
<output>
<ID>OUT</ID>520 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>676</ID>
<type>DA_FROM</type>
<position>-65.5,47</position>
<input>
<ID>IN_0</ID>523 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-STORE</lparam></gate>
<gate>
<ID>677</ID>
<type>DA_FROM</type>
<position>-66,38</position>
<input>
<ID>IN_0</ID>525 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-2</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>-43,40</position>
<input>
<ID>IN_0</ID>590 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE-RAM-WRITE</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>-51.5,44</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE-LOAD-MBR</lparam></gate>
<gate>
<ID>507</ID>
<type>DE_TO</type>
<position>-111.5,64.5</position>
<input>
<ID>IN_0</ID>565 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READ-SEQ-RESET</lparam></gate>
<gate>
<ID>121</ID>
<type>DE_TO</type>
<position>-116,9</position>
<input>
<ID>IN_0</ID>500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-MBR</lparam></gate>
<gate>
<ID>125</ID>
<type>DE_TO</type>
<position>-111.5,76.5</position>
<input>
<ID>IN_0</ID>379 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READ-LOAD-MBR</lparam></gate>
<gate>
<ID>324</ID>
<type>AA_LABEL</type>
<position>-61.5,52.5</position>
<gparam>LABEL_TEXT Store</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>325</ID>
<type>AA_LABEL</type>
<position>-89,-36.5</position>
<gparam>LABEL_TEXT Jump</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>715</ID>
<type>AA_LABEL</type>
<position>-123,18</position>
<gparam>LABEL_TEXT Add</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>716</ID>
<type>AA_LABEL</type>
<position>-59,20</position>
<gparam>LABEL_TEXT Sub</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>718</ID>
<type>DA_FROM</type>
<position>-65.5,43</position>
<input>
<ID>IN_0</ID>524 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-1</lparam></gate>
<gate>
<ID>719</ID>
<type>AA_AND2</type>
<position>-58,44</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>524 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>720</ID>
<type>AA_AND2</type>
<position>-58,39</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>525 </input>
<output>
<ID>OUT</ID>596 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>143</ID>
<type>DE_TO</type>
<position>-104,80.5</position>
<input>
<ID>IN_0</ID>381 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-IN</lparam></gate>
<gate>
<ID>339</ID>
<type>DE_TO</type>
<position>-40.5,-22.5</position>
<input>
<ID>IN_0</ID>513 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-R0</lparam></gate>
<gate>
<ID>340</ID>
<type>DE_TO</type>
<position>-40.5,-18</position>
<input>
<ID>IN_0</ID>509 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-R1</lparam></gate>
<gate>
<ID>341</ID>
<type>DA_FROM</type>
<position>-50.5,-14</position>
<input>
<ID>IN_0</ID>511 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID REG-SELECT</lparam></gate>
<gate>
<ID>342</ID>
<type>AA_AND2</type>
<position>-47,-18</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AE_OR2</type>
<position>-110.5,80.5</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>381 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>343</ID>
<type>AE_SMALL_INVERTER</type>
<position>-53,-18</position>
<input>
<ID>IN_0</ID>511 </input>
<output>
<ID>OUT_0</ID>514 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>344</ID>
<type>AA_AND2</type>
<position>-47,-22.5</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>512 </input>
<output>
<ID>OUT</ID>513 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>731</ID>
<type>DE_TO</type>
<position>-111.5,68</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READ-RAM-WRITE</lparam></gate>
<gate>
<ID>548</ID>
<type>AE_OR2</type>
<position>-109.5,72.5</position>
<input>
<ID>IN_0</ID>379 </input>
<input>
<ID>IN_1</ID>576 </input>
<output>
<ID>OUT</ID>575 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>552</ID>
<type>AE_OR2</type>
<position>-49.5,40</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>596 </input>
<output>
<ID>OUT</ID>590 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>553</ID>
<type>DA_FROM</type>
<position>-66,33</position>
<input>
<ID>IN_0</ID>589 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-3</lparam></gate>
<gate>
<ID>554</ID>
<type>AA_AND2</type>
<position>-58,34</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>589 </input>
<output>
<ID>OUT</ID>588 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>555</ID>
<type>DE_TO</type>
<position>-51.5,34</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE-SEQ-RESET</lparam></gate>
<gate>
<ID>749</ID>
<type>DE_TO</type>
<position>-116,-20</position>
<input>
<ID>IN_0</ID>462 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-SEQ-RESET</lparam></gate>
<gate>
<ID>750</ID>
<type>DE_TO</type>
<position>-52.5,-28</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-SEQ-RESET</lparam></gate>
<gate>
<ID>557</ID>
<type>DE_TO</type>
<position>-111.5,86.5</position>
<input>
<ID>IN_0</ID>483 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READ-PENDING</lparam></gate>
<gate>
<ID>751</ID>
<type>DA_FROM</type>
<position>-100.5,-43.5</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-JUMP</lparam></gate>
<gate>
<ID>1717</ID>
<type>AA_LABEL</type>
<position>-90,108</position>
<gparam>LABEL_TEXT Command Sequencing</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>559</ID>
<type>DE_TO</type>
<position>-54.5,80.5</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-OUT</lparam></gate>
<gate>
<ID>752</ID>
<type>DA_FROM</type>
<position>-101,-52.5</position>
<input>
<ID>IN_0</ID>571 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-2</lparam></gate>
<gate>
<ID>753</ID>
<type>DE_TO</type>
<position>-86.5,-51.5</position>
<input>
<ID>IN_0</ID>531 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JUMP-SEQ-RESET</lparam></gate>
<gate>
<ID>560</ID>
<type>DA_FROM</type>
<position>-68.5,88.5</position>
<input>
<ID>IN_0</ID>488 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OP-WRITE</lparam></gate>
<gate>
<ID>758</ID>
<type>DA_FROM</type>
<position>-100.5,-47.5</position>
<input>
<ID>IN_0</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-1</lparam></gate>
<gate>
<ID>760</ID>
<type>AA_AND2</type>
<position>-93,-46.5</position>
<input>
<ID>IN_0</ID>566 </input>
<input>
<ID>IN_1</ID>567 </input>
<output>
<ID>OUT</ID>585 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>761</ID>
<type>AA_AND2</type>
<position>-93,-51.5</position>
<input>
<ID>IN_0</ID>566 </input>
<input>
<ID>IN_1</ID>571 </input>
<output>
<ID>OUT</ID>531 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>DE_TO</type>
<position>-51.5,-9.5</position>
<input>
<ID>IN_0</ID>537 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-ADDER-RESULT</lparam></gate>
<gate>
<ID>575</ID>
<type>DA_FROM</type>
<position>-69,79.5</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-2</lparam></gate>
<gate>
<ID>382</ID>
<type>DE_TO</type>
<position>-52,-4.5</position>
<input>
<ID>IN_0</ID>540 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-ADDER</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>-69,74</position>
<input>
<ID>IN_0</ID>491 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-3</lparam></gate>
<gate>
<ID>577</ID>
<type>DA_FROM</type>
<position>-68.5,84.5</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-EXEC-1</lparam></gate>
<gate>
<ID>578</ID>
<type>AA_AND2</type>
<position>-61,85.5</position>
<input>
<ID>IN_0</ID>488 </input>
<input>
<ID>IN_1</ID>489 </input>
<output>
<ID>OUT</ID>492 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>584</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-82,-45.5,-80.5,-45.5</points>
<connection>
<GID>782</GID>
<name>IN_0</name></connection>
<intersection>-82 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-82,-45.5,-82,-45.5</points>
<connection>
<GID>774</GID>
<name>OUT</name></connection>
<intersection>-45.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>585</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,-46.5,-88,-46.5</points>
<connection>
<GID>760</GID>
<name>OUT</name></connection>
<connection>
<GID>774</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>588</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55,34,-53.5,34</points>
<connection>
<GID>555</GID>
<name>IN_0</name></connection>
<connection>
<GID>554</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>589</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-64,33,-61,33</points>
<connection>
<GID>554</GID>
<name>IN_1</name></connection>
<connection>
<GID>553</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>590</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46.5,40,-45,40</points>
<connection>
<GID>552</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>596</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-55,39,-52.5,39</points>
<connection>
<GID>552</GID>
<name>IN_1</name></connection>
<connection>
<GID>720</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,4,-118,4</points>
<connection>
<GID>663</GID>
<name>IN_0</name></connection>
<connection>
<GID>658</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,-1.5,-118,-1.5</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<connection>
<GID>659</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>608</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-28,-54.5,-28</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<connection>
<GID>652</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-67,69,-64,69</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<connection>
<GID>243</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,70,-56,70</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<connection>
<GID>243</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>636</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-83,-41.5,-80.5,-41.5</points>
<connection>
<GID>803</GID>
<name>IN_0</name></connection>
<connection>
<GID>778</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>637</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-88.5,-44.5,-88.5,-41.5</points>
<intersection>-44.5 1</intersection>
<intersection>-41.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-88.5,-44.5,-88,-44.5</points>
<connection>
<GID>774</GID>
<name>IN_0</name></connection>
<intersection>-88.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-88.5,-41.5,-87,-41.5</points>
<connection>
<GID>803</GID>
<name>OUT_0</name></connection>
<intersection>-88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120.5,29,-119,29</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>82</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-129.5,28,-126.5,28</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>451</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,80.5,-56.5,80.5</points>
<connection>
<GID>559</GID>
<name>IN_0</name></connection>
<connection>
<GID>613</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>452</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,75,-56.5,75</points>
<connection>
<GID>614</GID>
<name>OUT</name></connection>
<connection>
<GID>602</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>453</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120.5,46.5,-118.5,46.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<connection>
<GID>628</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,70.5,-121,70.5</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<connection>
<GID>84</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-107.5,-10.5,-106,-10.5</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<connection>
<GID>245</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116.5,-8.5,-113.5,-8.5</points>
<intersection>-116.5 44</intersection>
<intersection>-113.5 52</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>-116.5,-8.5,-116.5,-6.5</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>-8.5 1</intersection>
<intersection>-6.5 45</intersection></vsegment>
<hsegment>
<ID>45</ID>
<points>-116.5,-6.5,-116,-6.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>-116.5 44</intersection></hsegment>
<vsegment>
<ID>52</ID>
<points>-113.5,-9.5,-113.5,-8.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>-8.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>-118.5,-16,-113.5,-16</points>
<connection>
<GID>259</GID>
<name>IN_1</name></connection>
<intersection>-118.5 19</intersection>
<intersection>-115 22</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-118.5,-16,-118.5,-7</points>
<intersection>-16 11</intersection>
<intersection>-7 21</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>-120,-7,-118.5,-7</points>
<connection>
<GID>668</GID>
<name>OUT</name></connection>
<intersection>-118.5 19</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-115,-16,-115,-11.5</points>
<intersection>-16 11</intersection>
<intersection>-11.5 23</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>-115,-11.5,-113.5,-11.5</points>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>-115 22</intersection></hsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-107.5,-15,-106,-15</points>
<connection>
<GID>259</GID>
<name>OUT</name></connection>
<connection>
<GID>244</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>-116.5,-14,-116.5,-12.5</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>-14 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-116.5,-14,-113.5,-14</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>-116.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,-20,-118,-20</points>
<connection>
<GID>749</GID>
<name>IN_0</name></connection>
<connection>
<GID>670</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>464</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-27,-63,14</points>
<intersection>-27 13</intersection>
<intersection>-22.5 11</intersection>
<intersection>-8.5 9</intersection>
<intersection>-3.5 7</intersection>
<intersection>1.5 5</intersection>
<intersection>7 3</intersection>
<intersection>12 1</intersection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63,12,-61.5,12</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-64,14,-63,14</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-63,7,-61.5,7</points>
<connection>
<GID>647</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-63,1.5,-61.5,1.5</points>
<connection>
<GID>648</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-63,-3.5,-61.5,-3.5</points>
<connection>
<GID>649</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-63,-8.5,-61.5,-8.5</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-63,-22.5,-62,-22.5</points>
<connection>
<GID>651</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-63,-27,-62,-27</points>
<connection>
<GID>652</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>465</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-64,10,-61.5,10</points>
<connection>
<GID>646</GID>
<name>IN_1</name></connection>
<connection>
<GID>645</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>466</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-64.5,5,-61.5,5</points>
<connection>
<GID>647</GID>
<name>IN_1</name></connection>
<connection>
<GID>637</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>467</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-64.5,-0.5,-61.5,-0.5</points>
<connection>
<GID>648</GID>
<name>IN_1</name></connection>
<connection>
<GID>640</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>468</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-64.5,-5.5,-61.5,-5.5</points>
<connection>
<GID>649</GID>
<name>IN_1</name></connection>
<connection>
<GID>641</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>469</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-64.5,-10.5,-61.5,-10.5</points>
<connection>
<GID>650</GID>
<name>IN_1</name></connection>
<connection>
<GID>642</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>470</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-65,-24.5,-62,-24.5</points>
<connection>
<GID>651</GID>
<name>IN_1</name></connection>
<connection>
<GID>643</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>857</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,90,-104,90</points>
<connection>
<GID>1033</GID>
<name>OUT</name></connection>
<connection>
<GID>1031</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>471</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-65,-29,-62,-29</points>
<connection>
<GID>652</GID>
<name>IN_1</name></connection>
<connection>
<GID>644</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>858</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-113.5,91,-113.5,93.5</points>
<intersection>91 1</intersection>
<intersection>93.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-113.5,91,-112,91</points>
<connection>
<GID>1033</GID>
<name>IN_0</name></connection>
<intersection>-113.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-113.5,93.5,-109.5,93.5</points>
<connection>
<GID>1035</GID>
<name>IN_0</name></connection>
<intersection>-113.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>472</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-127.5,-19,-127.5,12</points>
<intersection>-19 17</intersection>
<intersection>-6 15</intersection>
<intersection>-0.5 5</intersection>
<intersection>5 3</intersection>
<intersection>10 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-127.5,10,-126,10</points>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>-127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-128.5,12,-127.5,12</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>-127.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-127.5,5,-126,5</points>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>-127.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-127.5,-0.5,-126,-0.5</points>
<connection>
<GID>659</GID>
<name>IN_0</name></connection>
<intersection>-127.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-127.5,-6,-126,-6</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<intersection>-127.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>-127.5,-19,-126,-19</points>
<connection>
<GID>670</GID>
<name>IN_0</name></connection>
<intersection>-127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>473</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-128.5,8,-126,8</points>
<connection>
<GID>657</GID>
<name>IN_1</name></connection>
<connection>
<GID>656</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>474</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-129,3,-126,3</points>
<connection>
<GID>658</GID>
<name>IN_1</name></connection>
<connection>
<GID>654</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>475</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-129,-2.5,-126,-2.5</points>
<connection>
<GID>659</GID>
<name>IN_1</name></connection>
<connection>
<GID>655</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>477</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-122.5,65.5,-122.5,89.5</points>
<intersection>65.5 18</intersection>
<intersection>72.5 12</intersection>
<intersection>77.5 5</intersection>
<intersection>82.5 3</intersection>
<intersection>87.5 1</intersection>
<intersection>89.5 10</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-122.5,87.5,-121,87.5</points>
<connection>
<GID>612</GID>
<name>IN_0</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-122.5,82.5,-121,82.5</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-122.5,77.5,-121,77.5</points>
<connection>
<GID>616</GID>
<name>IN_0</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-123.5,89.5,-122.5,89.5</points>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-122.5,72.5,-121,72.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>-122.5 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-122.5,65.5,-121,65.5</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>-122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>478</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-123.5,85.5,-121,85.5</points>
<connection>
<GID>612</GID>
<name>IN_1</name></connection>
<connection>
<GID>611</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>479</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,80.5,-121,80.5</points>
<connection>
<GID>615</GID>
<name>IN_1</name></connection>
<connection>
<GID>605</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>480</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-123.5,75.5,-121,75.5</points>
<connection>
<GID>616</GID>
<name>IN_1</name></connection>
<connection>
<GID>608</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>483</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115,86.5,-113.5,86.5</points>
<connection>
<GID>612</GID>
<name>OUT</name></connection>
<intersection>-113.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-113.5,86.5,-113.5,89</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<intersection>86.5 1</intersection>
<intersection>89 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-113.5,89,-112,89</points>
<connection>
<GID>1033</GID>
<name>IN_1</name></connection>
<intersection>-113.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>488</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65.5,71,-65.5,88.5</points>
<intersection>71 7</intersection>
<intersection>76 5</intersection>
<intersection>81.5 3</intersection>
<intersection>86.5 1</intersection>
<intersection>88.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65.5,86.5,-64,86.5</points>
<connection>
<GID>578</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66.5,88.5,-65.5,88.5</points>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-65.5,81.5,-64,81.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-65.5,76,-64,76</points>
<connection>
<GID>614</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-65.5,71,-64,71</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>-65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>489</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-66.5,84.5,-64,84.5</points>
<connection>
<GID>578</GID>
<name>IN_1</name></connection>
<connection>
<GID>577</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>490</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-67,79.5,-64,79.5</points>
<connection>
<GID>575</GID>
<name>IN_0</name></connection>
<connection>
<GID>613</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>491</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-67,74,-64,74</points>
<connection>
<GID>576</GID>
<name>IN_0</name></connection>
<connection>
<GID>614</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>492</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,85.5,-56.5,85.5</points>
<connection>
<GID>578</GID>
<name>OUT</name></connection>
<connection>
<GID>242</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>494</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-129,-8,-126,-8</points>
<connection>
<GID>669</GID>
<name>IN_0</name></connection>
<connection>
<GID>668</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>495</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-128,30,-128,49.5</points>
<intersection>30 5</intersection>
<intersection>42.5 3</intersection>
<intersection>47.5 1</intersection>
<intersection>49.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-128,47.5,-126.5,47.5</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-129,49.5,-128,49.5</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-128,42.5,-126.5,42.5</points>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-128,30,-126.5,30</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-128 0</intersection></hsegment></shape></wire>
<wire>
<ID>496</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-129,45.5,-126.5,45.5</points>
<connection>
<GID>628</GID>
<name>IN_1</name></connection>
<connection>
<GID>626</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>497</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-129.5,40.5,-126.5,40.5</points>
<connection>
<GID>631</GID>
<name>IN_1</name></connection>
<connection>
<GID>619</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>498</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-129,-21,-126,-21</points>
<connection>
<GID>671</GID>
<name>IN_0</name></connection>
<connection>
<GID>670</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>500</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120,9,-118,9</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>657</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>504</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55.5,11,-54,11</points>
<connection>
<GID>646</GID>
<name>OUT</name></connection>
<connection>
<GID>639</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>505</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55.5,6,-54,6</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<connection>
<GID>647</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>-55,44,-53.5,44</points>
<connection>
<GID>719</GID>
<name>OUT</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-53.5 19</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-53.5,41,-53.5,44</points>
<intersection>41 20</intersection>
<intersection>44 11</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-53.5,41,-52.5,41</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<intersection>-53.5 19</intersection></hsegment></shape></wire>
<wire>
<ID>509</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-44,-18,-42.5,-18</points>
<connection>
<GID>342</GID>
<name>OUT</name></connection>
<connection>
<GID>340</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>511</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-16,-50,-16</points>
<intersection>-53 44</intersection>
<intersection>-50 46</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>-53,-16,-53,-14</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>-16 1</intersection>
<intersection>-14 45</intersection></vsegment>
<hsegment>
<ID>45</ID>
<points>-53,-14,-52.5,-14</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<intersection>-53 44</intersection></hsegment>
<vsegment>
<ID>46</ID>
<points>-50,-17,-50,-16</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>512</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>-56,-23.5,-50,-23.5</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<connection>
<GID>651</GID>
<name>OUT</name></connection>
<intersection>-51.5 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>-51.5,-23.5,-51.5,-19</points>
<intersection>-23.5 11</intersection>
<intersection>-19 26</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>-51.5,-19,-50,-19</points>
<connection>
<GID>342</GID>
<name>IN_1</name></connection>
<intersection>-51.5 25</intersection></hsegment></shape></wire>
<wire>
<ID>513</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44,-22.5,-42.5,-22.5</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<connection>
<GID>339</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>514</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>-53,-21.5,-53,-20</points>
<connection>
<GID>343</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-53,-21.5,-50,-21.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>-53 6</intersection></hsegment></shape></wire>
<wire>
<ID>516</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-110,37.5,-108.5,37.5</points>
<connection>
<GID>672</GID>
<name>OUT</name></connection>
<connection>
<GID>662</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>517</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-119,39.5,-116,39.5</points>
<intersection>-119 44</intersection>
<intersection>-116 46</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>-119,39.5,-119,41.5</points>
<connection>
<GID>674</GID>
<name>IN_0</name></connection>
<intersection>39.5 1</intersection>
<intersection>41.5 45</intersection></vsegment>
<hsegment>
<ID>45</ID>
<points>-119,41.5,-118.5,41.5</points>
<connection>
<GID>666</GID>
<name>IN_0</name></connection>
<intersection>-119 44</intersection></hsegment>
<vsegment>
<ID>46</ID>
<points>-116,38.5,-116,39.5</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<intersection>39.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>518</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>-120.5,32,-116,32</points>
<connection>
<GID>675</GID>
<name>IN_1</name></connection>
<intersection>-120.5 19</intersection>
<intersection>-117.5 21</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>-120.5,32,-120.5,41.5</points>
<connection>
<GID>631</GID>
<name>OUT</name></connection>
<intersection>32 11</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>-117.5,32,-117.5,36.5</points>
<intersection>32 11</intersection>
<intersection>36.5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>-117.5,36.5,-116,36.5</points>
<connection>
<GID>672</GID>
<name>IN_1</name></connection>
<intersection>-117.5 21</intersection></hsegment></shape></wire>
<wire>
<ID>520</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-110,33,-108.5,33</points>
<connection>
<GID>675</GID>
<name>OUT</name></connection>
<connection>
<GID>661</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>521</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>-119,34,-119,35.5</points>
<connection>
<GID>674</GID>
<name>OUT_0</name></connection>
<intersection>34 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-119,34,-116,34</points>
<connection>
<GID>675</GID>
<name>IN_0</name></connection>
<intersection>-119 6</intersection></hsegment></shape></wire>
<wire>
<ID>523</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,35,-62.5,47</points>
<intersection>35 5</intersection>
<intersection>40 3</intersection>
<intersection>45 1</intersection>
<intersection>47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,45,-61,45</points>
<connection>
<GID>719</GID>
<name>IN_0</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63.5,47,-62.5,47</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-62.5,40,-61,40</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-62.5,35,-61,35</points>
<connection>
<GID>554</GID>
<name>IN_0</name></connection>
<intersection>-62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>524</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-63.5,43,-61,43</points>
<connection>
<GID>719</GID>
<name>IN_1</name></connection>
<connection>
<GID>718</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>525</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-64,38,-61,38</points>
<connection>
<GID>720</GID>
<name>IN_1</name></connection>
<connection>
<GID>677</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>531</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-90,-51.5,-88.5,-51.5</points>
<connection>
<GID>761</GID>
<name>OUT</name></connection>
<connection>
<GID>753</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>537</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55.5,-9.5,-53.5,-9.5</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<connection>
<GID>650</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>540</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55.5,-4.5,-54,-4.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<connection>
<GID>649</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>556</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55.5,0.5,-53.5,0.5</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<connection>
<GID>648</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>564</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,63.5,-121,63.5</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<connection>
<GID>459</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>565</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115,64.5,-113.5,64.5</points>
<connection>
<GID>507</GID>
<name>IN_0</name></connection>
<connection>
<GID>463</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>566</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-97.5,-50.5,-97.5,-43.5</points>
<intersection>-50.5 3</intersection>
<intersection>-45.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-97.5,-45.5,-96,-45.5</points>
<connection>
<GID>760</GID>
<name>IN_0</name></connection>
<intersection>-97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-98.5,-43.5,-97.5,-43.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<intersection>-97.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-97.5,-50.5,-96,-50.5</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<intersection>-97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>567</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-98.5,-47.5,-96,-47.5</points>
<connection>
<GID>760</GID>
<name>IN_1</name></connection>
<connection>
<GID>758</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>571</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-99,-52.5,-96,-52.5</points>
<connection>
<GID>761</GID>
<name>IN_1</name></connection>
<connection>
<GID>752</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>379</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-115,76.5,-115,79.5</points>
<connection>
<GID>616</GID>
<name>OUT</name></connection>
<intersection>76.5 13</intersection>
<intersection>79.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-115,79.5,-113.5,79.5</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-115 4</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-115,76.5,-113.5,76.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-115 4</intersection>
<intersection>-113.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-113.5,73.5,-113.5,76.5</points>
<intersection>73.5 15</intersection>
<intersection>76.5 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-113.5,73.5,-112.5,73.5</points>
<connection>
<GID>548</GID>
<name>IN_0</name></connection>
<intersection>-113.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>380</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-115,81.5,-113.5,81.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<connection>
<GID>615</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>381</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-107.5,80.5,-106,80.5</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<connection>
<GID>143</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>575</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-114,68,-114,69.5</points>
<intersection>68 3</intersection>
<intersection>69.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-114,69.5,-105.5,69.5</points>
<intersection>-114 0</intersection>
<intersection>-105.5 4</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-114,68,-113.5,68</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<intersection>-114 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-105.5,69.5,-105.5,72.5</points>
<intersection>69.5 2</intersection>
<intersection>72.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-106.5,72.5,-105.5,72.5</points>
<connection>
<GID>548</GID>
<name>OUT</name></connection>
<intersection>-105.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>576</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-115,71.5,-112.5,71.5</points>
<connection>
<GID>548</GID>
<name>IN_1</name></connection>
<connection>
<GID>86</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 7>
<page 8>
<PageViewport>-38.9938,296.788,182.618,184.766</PageViewport>
<gate>
<ID>772</ID>
<type>DA_FROM</type>
<position>52,251.5</position>
<input>
<ID>IN_0</ID>874 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-SEQ-RESET</lparam></gate>
<gate>
<ID>773</ID>
<type>DA_FROM</type>
<position>52,249.5</position>
<input>
<ID>IN_0</ID>873 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID JUMP-SEQ-RESET</lparam></gate>
<gate>
<ID>388</ID>
<type>AE_OR2</type>
<position>58,205</position>
<input>
<ID>IN_0</ID>455 </input>
<input>
<ID>IN_1</ID>456 </input>
<output>
<ID>OUT</ID>454 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>50.5,206</position>
<input>
<ID>IN_0</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-ADDER-RESULT</lparam></gate>
<gate>
<ID>783</ID>
<type>DA_FROM</type>
<position>51,224</position>
<input>
<ID>IN_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READ-RAM-WRITE</lparam></gate>
<gate>
<ID>785</ID>
<type>DA_FROM</type>
<position>51,222</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE-RAM-WRITE</lparam></gate>
<gate>
<ID>786</ID>
<type>DA_FROM</type>
<position>52,232</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-MBR</lparam></gate>
<gate>
<ID>788</ID>
<type>DE_TO</type>
<position>74,236</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-MBR</lparam></gate>
<gate>
<ID>793</ID>
<type>DA_FROM</type>
<position>52,230</position>
<input>
<ID>IN_0</ID>559 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READ-LOAD-MBR</lparam></gate>
<gate>
<ID>414</ID>
<type>DE_TO</type>
<position>65,205</position>
<input>
<ID>IN_0</ID>454 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-ADDER-RESULT</lparam></gate>
<gate>
<ID>416</ID>
<type>DA_FROM</type>
<position>50.5,204</position>
<input>
<ID>IN_0</ID>456 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-ADDER-RESULT</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_OR2</type>
<position>58,213.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>432</ID>
<type>AE_OR3</type>
<position>37.5,188</position>
<input>
<ID>IN_0</ID>486 </input>
<input>
<ID>IN_1</ID>487 </input>
<input>
<ID>IN_2</ID>476 </input>
<output>
<ID>OUT</ID>493 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>433</ID>
<type>AE_OR3</type>
<position>81.5,188</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>485 </input>
<input>
<ID>IN_2</ID>482 </input>
<output>
<ID>OUT</ID>499 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>434</ID>
<type>DA_FROM</type>
<position>75,188</position>
<input>
<ID>IN_0</ID>485 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-R1</lparam></gate>
<gate>
<ID>435</ID>
<type>DA_FROM</type>
<position>31,188</position>
<input>
<ID>IN_0</ID>487 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-R0</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>65.5,213.5</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-ADDER</lparam></gate>
<gate>
<ID>1020</ID>
<type>AE_OR2</type>
<position>58,197.5</position>
<input>
<ID>IN_0</ID>848 </input>
<input>
<ID>IN_1</ID>847 </input>
<output>
<ID>OUT</ID>849 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1021</ID>
<type>DA_FROM</type>
<position>50,198.5</position>
<input>
<ID>IN_0</ID>848 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLOCK-PULSE</lparam></gate>
<gate>
<ID>1022</ID>
<type>DA_FROM</type>
<position>50,196.5</position>
<input>
<ID>IN_0</ID>847 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PROGRAM-CLOCK-PULSE</lparam></gate>
<gate>
<ID>1023</ID>
<type>DE_TO</type>
<position>65,197.5</position>
<input>
<ID>IN_0</ID>849 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLOCK-PULSE-IN</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>55,268</position>
<gparam>LABEL_TEXT Conflict Resolution</gparam>
<gparam>TEXT_HEIGHT 1.4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>51.5,214.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-ADDER</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>51.5,212.5</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-ADDER</lparam></gate>
<gate>
<ID>68</ID>
<type>DA_FROM</type>
<position>52,239</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WRITE-LOAD-MBR</lparam></gate>
<gate>
<ID>74</ID>
<type>AE_OR3</type>
<position>58.5,232</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>559 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>77</ID>
<type>AE_OR2</type>
<position>66,236</position>
<input>
<ID>IN_0</ID>450 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1059</ID>
<type>AA_AND2</type>
<position>89,250.5</position>
<input>
<ID>IN_0</ID>507 </input>
<input>
<ID>IN_1</ID>872 </input>
<output>
<ID>OUT</ID>870 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1061</ID>
<type>DA_FROM</type>
<position>79,249.5</position>
<input>
<ID>IN_0</ID>871 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RESET-PC-IN</lparam></gate>
<gate>
<ID>1063</ID>
<type>AE_SMALL_INVERTER</type>
<position>83,249.5</position>
<input>
<ID>IN_0</ID>871 </input>
<output>
<ID>OUT_0</ID>872 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>1064</ID>
<type>DA_FROM</type>
<position>52,247.5</position>
<input>
<ID>IN_0</ID>876 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PROGRAM-SEQ-RESET</lparam></gate>
<gate>
<ID>1065</ID>
<type>AE_OR4</type>
<position>58.5,250.5</position>
<input>
<ID>IN_0</ID>875 </input>
<input>
<ID>IN_1</ID>874 </input>
<input>
<ID>IN_2</ID>873 </input>
<input>
<ID>IN_3</ID>876 </input>
<output>
<ID>OUT</ID>877 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>109</ID>
<type>DA_FROM</type>
<position>52,234</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE-LOAD-MBR</lparam></gate>
<gate>
<ID>887</ID>
<type>DE_TO</type>
<position>95.5,250.5</position>
<input>
<ID>IN_0</ID>870 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INCREMENT-PC</lparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>52,237</position>
<input>
<ID>IN_0</ID>580 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-LOAD-MBR</lparam></gate>
<gate>
<ID>326</ID>
<type>DA_FROM</type>
<position>52,241</position>
<input>
<ID>IN_0</ID>447 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-LOAD-MBR</lparam></gate>
<gate>
<ID>327</ID>
<type>DA_FROM</type>
<position>31,190</position>
<input>
<ID>IN_0</ID>486 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-LOAD-R0</lparam></gate>
<gate>
<ID>328</ID>
<type>DA_FROM</type>
<position>31,186</position>
<input>
<ID>IN_0</ID>476 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-R0</lparam></gate>
<gate>
<ID>330</ID>
<type>DE_TO</type>
<position>45,188</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-R0</lparam></gate>
<gate>
<ID>717</ID>
<type>DE_TO</type>
<position>73.5,255.5</position>
<input>
<ID>IN_0</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SEQ-RESET</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>75,190</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-LOAD-R1</lparam></gate>
<gate>
<ID>334</ID>
<type>DA_FROM</type>
<position>75,186</position>
<input>
<ID>IN_0</ID>482 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SUB-LOAD-R1</lparam></gate>
<gate>
<ID>335</ID>
<type>DE_TO</type>
<position>88,188</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-R1</lparam></gate>
<gate>
<ID>724</ID>
<type>AE_OR2</type>
<position>66.5,255.5</position>
<input>
<ID>IN_0</ID>532 </input>
<input>
<ID>IN_1</ID>877 </input>
<output>
<ID>OUT</ID>507 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>727</ID>
<type>AE_OR2</type>
<position>58,223</position>
<input>
<ID>IN_0</ID>562 </input>
<input>
<ID>IN_1</ID>563 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>728</ID>
<type>DE_TO</type>
<position>65,223</position>
<input>
<ID>IN_0</ID>510 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RAM-WRITE</lparam></gate>
<gate>
<ID>1718</ID>
<type>AA_LABEL</type>
<position>55.5,278</position>
<gparam>LABEL_TEXT Command Sequencing</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>755</ID>
<type>AE_OR4</type>
<position>58.5,259.5</position>
<input>
<ID>IN_0</ID>533 </input>
<input>
<ID>IN_1</ID>534 </input>
<input>
<ID>IN_2</ID>535 </input>
<input>
<ID>IN_3</ID>536 </input>
<output>
<ID>OUT</ID>532 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>757</ID>
<type>DA_FROM</type>
<position>52,262.5</position>
<input>
<ID>IN_0</ID>533 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID READ-SEQ-RESET</lparam></gate>
<gate>
<ID>763</ID>
<type>DA_FROM</type>
<position>52,260.5</position>
<input>
<ID>IN_0</ID>534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID WRITE-SEQ-RESET</lparam></gate>
<gate>
<ID>764</ID>
<type>DA_FROM</type>
<position>52,258.5</position>
<input>
<ID>IN_0</ID>535 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LOAD-SEQ-RESET</lparam></gate>
<gate>
<ID>383</ID>
<type>AE_OR3</type>
<position>58.5,239</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>448 </input>
<input>
<ID>IN_2</ID>580 </input>
<output>
<ID>OUT</ID>450 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>769</ID>
<type>DA_FROM</type>
<position>52,256.5</position>
<input>
<ID>IN_0</ID>536 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STORE-SEQ-RESET</lparam></gate>
<gate>
<ID>771</ID>
<type>DA_FROM</type>
<position>52,253.5</position>
<input>
<ID>IN_0</ID>875 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD-SEQ-RESET</lparam></gate>
<wire>
<ID>580</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,237,55.5,237</points>
<connection>
<GID>383</GID>
<name>IN_2</name></connection>
<connection>
<GID>124</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,213.5,63.5,213.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,214.5,55,214.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,212.5,55,212.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,232,55.5,232</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<connection>
<GID>786</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,234,55.5,234</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,232,62,235</points>
<intersection>232 3</intersection>
<intersection>235 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,235,63,235</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>61.5,232,62,232</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,236,72,236</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<connection>
<GID>788</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>447</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>54,241,55.5,241</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>448</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>54,239,55.5,239</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<connection>
<GID>68</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>450</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,237,62,239</points>
<intersection>237 4</intersection>
<intersection>239 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>61.5,239,62,239</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>62 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>62,237,63,237</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>62 0</intersection></hsegment></shape></wire>
<wire>
<ID>454</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,205,63,205</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<connection>
<GID>388</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>455</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,206,55,206</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<connection>
<GID>388</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52.5,204,55,204</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<connection>
<GID>388</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>847</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,196.5,55,196.5</points>
<connection>
<GID>1022</GID>
<name>IN_0</name></connection>
<connection>
<GID>1020</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>848</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>52,198.5,55,198.5</points>
<connection>
<GID>1021</GID>
<name>IN_0</name></connection>
<connection>
<GID>1020</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>849</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>61,197.5,63,197.5</points>
<connection>
<GID>1023</GID>
<name>IN_0</name></connection>
<connection>
<GID>1020</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>476</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>33,186,34.5,186</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<connection>
<GID>432</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>482</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>77,186,78.5,186</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>870</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92,250.5,93.5,250.5</points>
<connection>
<GID>887</GID>
<name>IN_0</name></connection>
<connection>
<GID>1059</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>484</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,190,78.5,190</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>871</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>81,249.5,81,249.5</points>
<connection>
<GID>1063</GID>
<name>IN_0</name></connection>
<connection>
<GID>1061</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>485</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,188,78.5,188</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>872</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>85,249.5,86,249.5</points>
<connection>
<GID>1059</GID>
<name>IN_1</name></connection>
<connection>
<GID>1063</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>486</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,190,34.5,190</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<connection>
<GID>432</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>873</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,249.5,55.5,249.5</points>
<connection>
<GID>773</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>487</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,188,34.5,188</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<connection>
<GID>432</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>874</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,251.5,55.5,251.5</points>
<connection>
<GID>772</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>875</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,253.5,55.5,253.5</points>
<connection>
<GID>771</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>876</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,247.5,55.5,247.5</points>
<connection>
<GID>1064</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>877</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,250.5,63,254.5</points>
<intersection>250.5 3</intersection>
<intersection>254.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>63,254.5,63.5,254.5</points>
<connection>
<GID>724</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>62.5,250.5,63,250.5</points>
<connection>
<GID>1065</GID>
<name>OUT</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>493</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40.5,188,43,188</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<connection>
<GID>432</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>499</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>84.5,188,86,188</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>507</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,255.5,71.5,255.5</points>
<connection>
<GID>717</GID>
<name>IN_0</name></connection>
<connection>
<GID>724</GID>
<name>OUT</name></connection>
<intersection>71.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>71.5,251.5,71.5,255.5</points>
<intersection>251.5 7</intersection>
<intersection>255.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>71.5,251.5,86,251.5</points>
<connection>
<GID>1059</GID>
<name>IN_0</name></connection>
<intersection>71.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>510</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>61,223,63,223</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<connection>
<GID>727</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>532</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,256.5,63,259.5</points>
<intersection>256.5 4</intersection>
<intersection>259.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62.5,259.5,63,259.5</points>
<connection>
<GID>755</GID>
<name>OUT</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>63,256.5,63.5,256.5</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>533</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,262.5,55.5,262.5</points>
<connection>
<GID>757</GID>
<name>IN_0</name></connection>
<connection>
<GID>755</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>534</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,260.5,55.5,260.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<connection>
<GID>755</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>535</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,258.5,55.5,258.5</points>
<connection>
<GID>764</GID>
<name>IN_0</name></connection>
<connection>
<GID>755</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>536</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,256.5,55.5,256.5</points>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<connection>
<GID>755</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>559</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,230,55.5,230</points>
<connection>
<GID>74</GID>
<name>IN_2</name></connection>
<connection>
<GID>793</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>562</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,224,55,224</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<connection>
<GID>783</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>563</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,222,55,222</points>
<connection>
<GID>727</GID>
<name>IN_1</name></connection>
<connection>
<GID>785</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>-56.9809,18.0487,64.3821,-43.2987</PageViewport>
<gate>
<ID>982</ID>
<type>AE_OR4</type>
<position>-16.5,-15</position>
<input>
<ID>IN_0</ID>819 </input>
<input>
<ID>IN_1</ID>821 </input>
<input>
<ID>IN_2</ID>820 </input>
<input>
<ID>IN_3</ID>818 </input>
<output>
<ID>OUT</ID>822 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>998</ID>
<type>BB_CLOCK</type>
<position>-12,2</position>
<output>
<ID>CLK</ID>856 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 10</lparam></gate>
<gate>
<ID>1000</ID>
<type>DE_TO</type>
<position>6.5,-4.5</position>
<input>
<ID>IN_0</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PROGRAM-CLOCK-PULSE</lparam></gate>
<gate>
<ID>816</ID>
<type>AA_LABEL</type>
<position>-4.5,8.5</position>
<gparam>LABEL_TEXT Program</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>823</ID>
<type>DA_FROM</type>
<position>-15.5,-9</position>
<input>
<ID>IN_0</ID>786 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RUN-PROGRAM</lparam></gate>
<gate>
<ID>1025</ID>
<type>AA_AND3</type>
<position>0.5,-4.5</position>
<input>
<ID>IN_0</ID>856 </input>
<input>
<ID>IN_1</ID>860 </input>
<input>
<ID>IN_2</ID>786 </input>
<output>
<ID>OUT</ID>851 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1027</ID>
<type>DA_FROM</type>
<position>-20,-5.5</position>
<input>
<ID>IN_0</ID>854 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID STOP-EXECUTION</lparam></gate>
<gate>
<ID>1029</ID>
<type>AE_SMALL_INVERTER</type>
<position>-15,-5.5</position>
<input>
<ID>IN_0</ID>854 </input>
<output>
<ID>OUT_0</ID>861 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>846</ID>
<type>DE_TO</type>
<position>12.5,-23</position>
<input>
<ID>IN_0</ID>686 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RESET-PC-IN</lparam></gate>
<gate>
<ID>1041</ID>
<type>DA_FROM</type>
<position>-15.5,-2</position>
<input>
<ID>IN_0</ID>862 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CONTINUE-PROGRAM</lparam></gate>
<gate>
<ID>849</ID>
<type>DA_FROM</type>
<position>-0.5,-24</position>
<input>
<ID>IN_0</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID RESET-PC</lparam></gate>
<gate>
<ID>1044</ID>
<type>AE_OR2</type>
<position>-8.5,-4.5</position>
<input>
<ID>IN_0</ID>862 </input>
<input>
<ID>IN_1</ID>861 </input>
<output>
<ID>OUT</ID>860 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>851</ID>
<type>AE_OR2</type>
<position>6,-23</position>
<input>
<ID>IN_0</ID>787 </input>
<input>
<ID>IN_1</ID>643 </input>
<output>
<ID>OUT</ID>686 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>856</ID>
<type>DA_FROM</type>
<position>-23,-14</position>
<input>
<ID>IN_0</ID>821 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-2</lparam></gate>
<gate>
<ID>859</ID>
<type>DA_FROM</type>
<position>-23,-18</position>
<input>
<ID>IN_0</ID>818 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-0</lparam></gate>
<gate>
<ID>871</ID>
<type>DA_FROM</type>
<position>-23,-12</position>
<input>
<ID>IN_0</ID>819 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-3</lparam></gate>
<gate>
<ID>1069</ID>
<type>DE_TO</type>
<position>12.5,-25</position>
<input>
<ID>IN_0</ID>686 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PROGRAM-SEQ-RESET</lparam></gate>
<gate>
<ID>890</ID>
<type>DA_FROM</type>
<position>-23,-16</position>
<input>
<ID>IN_0</ID>820 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC-1</lparam></gate>
<gate>
<ID>950</ID>
<type>DA_FROM</type>
<position>-23,-20.5</position>
<input>
<ID>IN_0</ID>782 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-REG-IN</lparam></gate>
<gate>
<ID>951</ID>
<type>DA_FROM</type>
<position>-23,-22.5</position>
<input>
<ID>IN_0</ID>783 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-3-IN</lparam></gate>
<gate>
<ID>952</ID>
<type>DA_FROM</type>
<position>-23,-24.5</position>
<input>
<ID>IN_0</ID>781 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-2-IN</lparam></gate>
<gate>
<ID>953</ID>
<type>DA_FROM</type>
<position>-23,-26.5</position>
<input>
<ID>IN_0</ID>780 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-1-IN</lparam></gate>
<gate>
<ID>954</ID>
<type>DA_FROM</type>
<position>-23,-28.5</position>
<input>
<ID>IN_0</ID>779 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-ADDR-0-IN</lparam></gate>
<gate>
<ID>955</ID>
<type>DA_FROM</type>
<position>-23,-30.5</position>
<input>
<ID>IN_0</ID>778 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-2-IN</lparam></gate>
<gate>
<ID>956</ID>
<type>DA_FROM</type>
<position>-23,-32.5</position>
<input>
<ID>IN_0</ID>777 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-1-IN</lparam></gate>
<gate>
<ID>957</ID>
<type>DA_FROM</type>
<position>-23,-34.5</position>
<input>
<ID>IN_0</ID>776 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR-OP-0-IN</lparam></gate>
<gate>
<ID>958</ID>
<type>DM_NOR8</type>
<position>-16.5,-27.5</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>783 </input>
<input>
<ID>IN_2</ID>781 </input>
<input>
<ID>IN_3</ID>780 </input>
<input>
<ID>IN_4</ID>776 </input>
<input>
<ID>IN_5</ID>777 </input>
<input>
<ID>IN_6</ID>778 </input>
<input>
<ID>IN_7</ID>779 </input>
<output>
<ID>OUT</ID>784 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>960</ID>
<type>AA_AND3</type>
<position>-7.5,-18.5</position>
<input>
<ID>IN_0</ID>786 </input>
<input>
<ID>IN_1</ID>822 </input>
<input>
<ID>IN_2</ID>784 </input>
<output>
<ID>OUT</ID>787 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<wire>
<ID>776</ID>
<shape>
<vsegment>
<ID>10</ID>
<points>-19.5,-34.5,-19.5,-31</points>
<connection>
<GID>958</GID>
<name>IN_4</name></connection>
<intersection>-34.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-21,-34.5,-19.5,-34.5</points>
<connection>
<GID>957</GID>
<name>IN_0</name></connection>
<intersection>-19.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>777</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-32.5,-20,-30</points>
<intersection>-32.5 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-20,-30,-19.5,-30</points>
<connection>
<GID>958</GID>
<name>IN_5</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-21,-32.5,-20,-32.5</points>
<connection>
<GID>956</GID>
<name>IN_0</name></connection>
<intersection>-20 0</intersection></hsegment></shape></wire>
<wire>
<ID>778</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-30.5,-20.5,-29</points>
<intersection>-30.5 8</intersection>
<intersection>-29 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-20.5,-29,-19.5,-29</points>
<connection>
<GID>958</GID>
<name>IN_6</name></connection>
<intersection>-20.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-21,-30.5,-20.5,-30.5</points>
<connection>
<GID>955</GID>
<name>IN_0</name></connection>
<intersection>-20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>779</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-28.5,-19.5,-28.5</points>
<connection>
<GID>954</GID>
<name>IN_0</name></connection>
<intersection>-19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19.5,-28.5,-19.5,-28</points>
<connection>
<GID>958</GID>
<name>IN_7</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>780</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-26.5,-19.5,-26.5</points>
<connection>
<GID>953</GID>
<name>IN_0</name></connection>
<intersection>-19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19.5,-27,-19.5,-26.5</points>
<connection>
<GID>958</GID>
<name>IN_3</name></connection>
<intersection>-26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>781</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-26,-20.5,-24.5</points>
<intersection>-26 2</intersection>
<intersection>-24.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-20.5,-26,-19.5,-26</points>
<connection>
<GID>958</GID>
<name>IN_2</name></connection>
<intersection>-20.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-21,-24.5,-20.5,-24.5</points>
<connection>
<GID>952</GID>
<name>IN_0</name></connection>
<intersection>-20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>782</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-24,-19.5,-20.5</points>
<connection>
<GID>958</GID>
<name>IN_0</name></connection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-20.5,-19.5,-20.5</points>
<connection>
<GID>950</GID>
<name>IN_0</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>783</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-25,-20,-22.5</points>
<intersection>-25 3</intersection>
<intersection>-22.5 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-20,-25,-19.5,-25</points>
<connection>
<GID>958</GID>
<name>IN_1</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-21,-22.5,-20,-22.5</points>
<connection>
<GID>951</GID>
<name>IN_0</name></connection>
<intersection>-20 0</intersection></hsegment></shape></wire>
<wire>
<ID>784</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-27.5,-12,-20.5</points>
<intersection>-27.5 5</intersection>
<intersection>-20.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-12,-20.5,-10.5,-20.5</points>
<connection>
<GID>960</GID>
<name>IN_2</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-12.5,-27.5,-12,-27.5</points>
<connection>
<GID>958</GID>
<name>OUT</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>786</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-9,-4,-9</points>
<connection>
<GID>823</GID>
<name>IN_0</name></connection>
<intersection>-11.5 26</intersection>
<intersection>-4 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>-4,-9,-4,-6.5</points>
<intersection>-9 1</intersection>
<intersection>-6.5 23</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>-4,-6.5,-2.5,-6.5</points>
<connection>
<GID>1025</GID>
<name>IN_2</name></connection>
<intersection>-4 22</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>-11.5,-16.5,-11.5,-9</points>
<intersection>-16.5 27</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>-11.5,-16.5,-10.5,-16.5</points>
<connection>
<GID>960</GID>
<name>IN_0</name></connection>
<intersection>-11.5 26</intersection></hsegment></shape></wire>
<wire>
<ID>787</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-22,-0.5,-18.5</points>
<intersection>-22 6</intersection>
<intersection>-18.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-4.5,-18.5,-0.5,-18.5</points>
<connection>
<GID>960</GID>
<name>OUT</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-0.5,-22,3,-22</points>
<connection>
<GID>851</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>818</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-18,-19.5,-18</points>
<connection>
<GID>982</GID>
<name>IN_3</name></connection>
<connection>
<GID>859</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>819</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-12,-19.5,-12</points>
<connection>
<GID>982</GID>
<name>IN_0</name></connection>
<connection>
<GID>871</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>820</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-16,-19.5,-16</points>
<connection>
<GID>982</GID>
<name>IN_2</name></connection>
<connection>
<GID>890</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>821</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-14,-19.5,-14</points>
<connection>
<GID>982</GID>
<name>IN_1</name></connection>
<connection>
<GID>856</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>822</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-18.5,-12.5,-15</points>
<connection>
<GID>982</GID>
<name>OUT</name></connection>
<intersection>-18.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-12.5,-18.5,-10.5,-18.5</points>
<connection>
<GID>960</GID>
<name>IN_1</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>643</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>1.5,-24,3,-24</points>
<connection>
<GID>849</GID>
<name>IN_0</name></connection>
<connection>
<GID>851</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>851</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-4.5,4.5,-4.5</points>
<connection>
<GID>1025</GID>
<name>OUT</name></connection>
<connection>
<GID>1000</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>854</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-18,-5.5,-17,-5.5</points>
<connection>
<GID>1027</GID>
<name>IN_0</name></connection>
<connection>
<GID>1029</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>856</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-2.5,-4,2</points>
<intersection>-2.5 3</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-8,2,-4,2</points>
<connection>
<GID>998</GID>
<name>CLK</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4,-2.5,-2.5,-2.5</points>
<connection>
<GID>1025</GID>
<name>IN_0</name></connection>
<intersection>-4 0</intersection></hsegment></shape></wire>
<wire>
<ID>860</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-5.5,-4.5,-2.5,-4.5</points>
<connection>
<GID>1025</GID>
<name>IN_1</name></connection>
<connection>
<GID>1044</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>861</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,-5.5,-11.5,-5.5</points>
<connection>
<GID>1044</GID>
<name>IN_1</name></connection>
<connection>
<GID>1029</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>862</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,-2,-11.5,-2</points>
<connection>
<GID>1041</GID>
<name>IN_0</name></connection>
<intersection>-11.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-11.5,-3.5,-11.5,-2</points>
<connection>
<GID>1044</GID>
<name>IN_0</name></connection>
<intersection>-2 1</intersection></vsegment></shape></wire>
<wire>
<ID>686</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>9,-23,10.5,-23</points>
<connection>
<GID>851</GID>
<name>OUT</name></connection>
<connection>
<GID>846</GID>
<name>IN_0</name></connection>
<intersection>10.5 29</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>10.5,-25,10.5,-23</points>
<connection>
<GID>1069</GID>
<name>IN_0</name></connection>
<intersection>-23 0</intersection></vsegment></shape></wire></page 9></circuit>